magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1510 582
<< pwell >>
rect 1 21 1471 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 247 47 277 177
rect 331 47 361 177
rect 415 47 445 177
rect 499 47 529 177
rect 583 47 613 177
rect 667 47 697 177
rect 751 47 781 177
rect 848 47 878 177
rect 934 47 964 177
rect 1019 47 1049 177
rect 1103 47 1133 177
rect 1187 47 1217 177
rect 1271 47 1301 177
rect 1357 47 1387 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 331 297 361 497
rect 415 297 445 497
rect 499 297 529 497
rect 583 297 613 497
rect 667 297 697 497
rect 751 297 781 497
rect 835 297 865 497
rect 919 297 949 497
rect 1009 297 1039 497
rect 1095 297 1125 497
rect 1181 297 1211 497
rect 1271 297 1301 497
rect 1363 297 1393 497
<< ndiff >>
rect 27 93 79 177
rect 27 59 35 93
rect 69 59 79 93
rect 27 47 79 59
rect 109 157 163 177
rect 109 123 119 157
rect 153 123 163 157
rect 109 47 163 123
rect 193 89 247 177
rect 193 55 203 89
rect 237 55 247 89
rect 193 47 247 55
rect 277 89 331 177
rect 277 55 287 89
rect 321 55 331 89
rect 277 47 331 55
rect 361 169 415 177
rect 361 135 371 169
rect 405 135 415 169
rect 361 47 415 135
rect 445 89 499 177
rect 445 55 455 89
rect 489 55 499 89
rect 445 47 499 55
rect 529 169 583 177
rect 529 135 539 169
rect 573 135 583 169
rect 529 47 583 135
rect 613 89 667 177
rect 613 55 623 89
rect 657 55 667 89
rect 613 47 667 55
rect 697 89 751 177
rect 697 55 707 89
rect 741 55 751 89
rect 697 47 751 55
rect 781 169 848 177
rect 781 135 795 169
rect 829 135 848 169
rect 781 101 848 135
rect 781 67 795 101
rect 829 67 848 101
rect 781 47 848 67
rect 878 89 934 177
rect 878 55 889 89
rect 923 55 934 89
rect 878 47 934 55
rect 964 169 1019 177
rect 964 135 975 169
rect 1009 135 1019 169
rect 964 101 1019 135
rect 964 67 975 101
rect 1009 67 1019 101
rect 964 47 1019 67
rect 1049 89 1103 177
rect 1049 55 1059 89
rect 1093 55 1103 89
rect 1049 47 1103 55
rect 1133 169 1187 177
rect 1133 135 1143 169
rect 1177 135 1187 169
rect 1133 101 1187 135
rect 1133 67 1143 101
rect 1177 67 1187 101
rect 1133 47 1187 67
rect 1217 89 1271 177
rect 1217 55 1227 89
rect 1261 55 1271 89
rect 1217 47 1271 55
rect 1301 165 1357 177
rect 1301 131 1313 165
rect 1347 131 1357 165
rect 1301 47 1357 131
rect 1387 89 1445 177
rect 1387 55 1399 89
rect 1433 55 1445 89
rect 1387 47 1445 55
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 297 79 375
rect 109 485 163 497
rect 109 451 119 485
rect 153 451 163 485
rect 109 297 163 451
rect 193 477 247 497
rect 193 443 203 477
rect 237 443 247 477
rect 193 409 247 443
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 489 331 497
rect 277 455 287 489
rect 321 455 331 489
rect 277 297 331 455
rect 361 477 415 497
rect 361 443 371 477
rect 405 443 415 477
rect 361 409 415 443
rect 361 375 371 409
rect 405 375 415 409
rect 361 297 415 375
rect 445 489 499 497
rect 445 455 455 489
rect 489 455 499 489
rect 445 297 499 455
rect 529 477 583 497
rect 529 443 539 477
rect 573 443 583 477
rect 529 409 583 443
rect 529 375 539 409
rect 573 375 583 409
rect 529 297 583 375
rect 613 489 667 497
rect 613 455 623 489
rect 657 455 667 489
rect 613 297 667 455
rect 697 477 751 497
rect 697 443 707 477
rect 741 443 751 477
rect 697 409 751 443
rect 697 375 707 409
rect 741 375 751 409
rect 697 297 751 375
rect 781 417 835 497
rect 781 383 791 417
rect 825 383 835 417
rect 781 297 835 383
rect 865 489 919 497
rect 865 455 875 489
rect 909 455 919 489
rect 865 297 919 455
rect 949 297 1009 497
rect 1039 413 1095 497
rect 1039 379 1050 413
rect 1084 379 1095 413
rect 1039 297 1095 379
rect 1125 339 1181 497
rect 1125 305 1136 339
rect 1170 305 1181 339
rect 1125 297 1181 305
rect 1211 413 1271 497
rect 1211 379 1226 413
rect 1260 379 1271 413
rect 1211 297 1271 379
rect 1301 297 1363 497
rect 1393 485 1445 497
rect 1393 451 1403 485
rect 1437 451 1445 485
rect 1393 297 1445 451
<< ndiffc >>
rect 35 59 69 93
rect 119 123 153 157
rect 203 55 237 89
rect 287 55 321 89
rect 371 135 405 169
rect 455 55 489 89
rect 539 135 573 169
rect 623 55 657 89
rect 707 55 741 89
rect 795 135 829 169
rect 795 67 829 101
rect 889 55 923 89
rect 975 135 1009 169
rect 975 67 1009 101
rect 1059 55 1093 89
rect 1143 135 1177 169
rect 1143 67 1177 101
rect 1227 55 1261 89
rect 1313 131 1347 165
rect 1399 55 1433 89
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 451 153 485
rect 203 443 237 477
rect 203 375 237 409
rect 287 455 321 489
rect 371 443 405 477
rect 371 375 405 409
rect 455 455 489 489
rect 539 443 573 477
rect 539 375 573 409
rect 623 455 657 489
rect 707 443 741 477
rect 707 375 741 409
rect 791 383 825 417
rect 875 455 909 489
rect 1050 379 1084 413
rect 1136 305 1170 339
rect 1226 379 1260 413
rect 1403 451 1437 485
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 331 497 361 523
rect 415 497 445 523
rect 499 497 529 523
rect 583 497 613 523
rect 667 497 697 523
rect 751 497 781 523
rect 835 497 865 523
rect 919 497 949 523
rect 1009 497 1039 523
rect 1095 497 1125 523
rect 1181 497 1211 523
rect 1271 497 1301 523
rect 1363 497 1393 523
rect 79 259 109 297
rect 163 259 193 297
rect 247 259 277 297
rect 75 249 277 259
rect 75 215 91 249
rect 125 215 159 249
rect 193 215 227 249
rect 261 215 277 249
rect 75 205 277 215
rect 79 177 109 205
rect 163 177 193 205
rect 247 177 277 205
rect 331 259 361 297
rect 415 259 445 297
rect 499 259 529 297
rect 583 259 613 297
rect 667 265 697 297
rect 751 265 781 297
rect 835 265 865 297
rect 919 265 949 297
rect 1009 265 1039 297
rect 1095 265 1125 297
rect 1181 265 1211 297
rect 1271 265 1301 297
rect 1363 265 1393 297
rect 331 249 613 259
rect 331 215 347 249
rect 381 215 415 249
rect 449 215 483 249
rect 517 215 551 249
rect 585 215 613 249
rect 331 205 613 215
rect 331 177 361 205
rect 415 177 445 205
rect 499 177 529 205
rect 583 177 613 205
rect 655 249 709 265
rect 655 215 665 249
rect 699 215 709 249
rect 655 199 709 215
rect 751 249 964 265
rect 751 215 765 249
rect 799 215 833 249
rect 867 215 901 249
rect 935 215 964 249
rect 751 199 964 215
rect 1006 249 1301 265
rect 1006 215 1016 249
rect 1050 215 1084 249
rect 1118 215 1152 249
rect 1186 215 1220 249
rect 1254 215 1301 249
rect 1006 199 1301 215
rect 1343 249 1398 265
rect 1343 215 1353 249
rect 1387 215 1398 249
rect 1343 199 1398 215
rect 667 177 697 199
rect 751 177 781 199
rect 848 177 878 199
rect 934 177 964 199
rect 1019 177 1049 199
rect 1103 177 1133 199
rect 1187 177 1217 199
rect 1271 177 1301 199
rect 1357 177 1387 199
rect 79 21 109 47
rect 163 21 193 47
rect 247 21 277 47
rect 331 21 361 47
rect 415 21 445 47
rect 499 21 529 47
rect 583 21 613 47
rect 667 21 697 47
rect 751 21 781 47
rect 848 21 878 47
rect 934 21 964 47
rect 1019 21 1049 47
rect 1103 21 1133 47
rect 1187 21 1217 47
rect 1271 21 1301 47
rect 1357 21 1387 47
<< polycont >>
rect 91 215 125 249
rect 159 215 193 249
rect 227 215 261 249
rect 347 215 381 249
rect 415 215 449 249
rect 483 215 517 249
rect 551 215 585 249
rect 665 215 699 249
rect 765 215 799 249
rect 833 215 867 249
rect 901 215 935 249
rect 1016 215 1050 249
rect 1084 215 1118 249
rect 1152 215 1186 249
rect 1220 215 1254 249
rect 1353 215 1387 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 19 477 69 493
rect 19 443 35 477
rect 103 485 169 527
rect 103 451 119 485
rect 153 451 169 485
rect 203 477 237 493
rect 19 417 69 443
rect 271 489 337 527
rect 271 455 287 489
rect 321 455 337 489
rect 371 477 405 493
rect 203 421 237 443
rect 439 489 505 527
rect 439 455 455 489
rect 489 455 505 489
rect 539 477 573 493
rect 371 421 405 443
rect 607 489 673 527
rect 607 455 623 489
rect 657 455 673 489
rect 707 489 1454 493
rect 707 477 875 489
rect 539 421 573 443
rect 741 455 875 477
rect 909 485 1454 489
rect 909 455 1403 485
rect 741 451 1403 455
rect 1437 451 1454 485
rect 707 421 741 443
rect 203 417 741 421
rect 19 409 741 417
rect 19 375 35 409
rect 69 375 203 409
rect 237 375 371 409
rect 405 375 539 409
rect 573 375 707 409
rect 19 359 741 375
rect 775 383 791 417
rect 825 383 982 417
rect 775 357 982 383
rect 1034 413 1455 417
rect 1034 379 1050 413
rect 1084 379 1226 413
rect 1260 379 1455 413
rect 1034 373 1455 379
rect 926 339 982 357
rect 20 289 715 325
rect 20 249 277 289
rect 332 249 601 255
rect 20 215 91 249
rect 125 215 159 249
rect 193 215 227 249
rect 261 215 277 249
rect 331 215 347 249
rect 381 215 415 249
rect 449 215 483 249
rect 517 215 551 249
rect 585 215 601 249
rect 20 207 277 215
rect 332 207 601 215
rect 649 249 715 289
rect 649 215 665 249
rect 699 215 715 249
rect 649 207 715 215
rect 749 289 766 323
rect 800 289 892 323
rect 926 305 1136 339
rect 1170 305 1192 339
rect 926 289 1192 305
rect 749 255 892 289
rect 1226 255 1270 339
rect 749 249 951 255
rect 749 215 765 249
rect 799 215 833 249
rect 867 215 901 249
rect 935 215 951 249
rect 749 207 951 215
rect 1000 249 1270 255
rect 1000 215 1016 249
rect 1050 215 1084 249
rect 1118 215 1152 249
rect 1186 215 1220 249
rect 1254 215 1270 249
rect 1000 207 1270 215
rect 1386 299 1455 373
rect 1318 265 1352 289
rect 1318 249 1387 265
rect 1318 215 1353 249
rect 1318 199 1387 215
rect 113 157 321 173
rect 113 123 119 157
rect 153 139 321 157
rect 153 123 155 139
rect 19 93 79 117
rect 113 106 155 123
rect 19 59 35 93
rect 69 59 79 93
rect 19 17 79 59
rect 190 89 237 105
rect 190 55 203 89
rect 190 17 237 55
rect 271 101 321 139
rect 355 169 1271 173
rect 355 135 371 169
rect 405 135 539 169
rect 573 139 795 169
rect 573 135 666 139
rect 775 135 795 139
rect 829 135 975 169
rect 1009 135 1143 169
rect 1177 165 1271 169
rect 1421 165 1455 299
rect 1177 135 1313 165
rect 775 131 1313 135
rect 1347 131 1455 165
rect 775 125 1455 131
rect 775 123 1009 125
rect 271 89 673 101
rect 271 55 287 89
rect 321 55 455 89
rect 489 55 623 89
rect 657 55 673 89
rect 271 51 673 55
rect 707 89 741 105
rect 707 17 741 55
rect 775 101 839 123
rect 775 67 795 101
rect 829 67 839 101
rect 975 101 1009 123
rect 775 51 839 67
rect 873 55 889 89
rect 923 55 939 89
rect 873 17 939 55
rect 1143 123 1455 125
rect 1143 101 1177 123
rect 975 51 1009 67
rect 1043 55 1059 89
rect 1093 55 1109 89
rect 1043 17 1109 55
rect 1143 51 1177 67
rect 1211 55 1227 89
rect 1261 55 1277 89
rect 1211 17 1277 55
rect 1383 55 1399 89
rect 1433 55 1454 89
rect 1383 17 1454 55
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 766 289 800 323
rect 1318 289 1352 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
<< metal1 >>
rect 0 561 1472 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1472 561
rect 0 496 1472 527
rect 754 323 812 329
rect 754 289 766 323
rect 800 320 812 323
rect 1306 323 1364 329
rect 1306 320 1318 323
rect 800 292 1318 320
rect 800 289 812 292
rect 754 283 812 289
rect 1306 289 1318 292
rect 1352 289 1364 323
rect 1306 283 1364 289
rect 0 17 1472 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1472 17
rect 0 -48 1472 -17
<< labels >>
flabel locali s 214 289 248 323 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 398 221 432 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 1042 221 1076 255 0 FreeSans 340 0 0 0 C1
port 4 nsew signal input
flabel locali s 1410 357 1444 391 0 FreeSans 340 0 0 0 Y
port 9 nsew signal output
flabel metal1 s 766 289 800 323 0 FreeSans 400 0 0 0 B1
port 3 nsew signal input
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
rlabel comment s 0 0 0 0 4 a211oi_4
rlabel locali s 1318 265 1352 323 1 B1
port 3 nsew signal input
rlabel locali s 1318 199 1387 265 1 B1
port 3 nsew signal input
rlabel metal1 s 1306 320 1364 329 1 B1
port 3 nsew signal input
rlabel metal1 s 1306 283 1364 292 1 B1
port 3 nsew signal input
rlabel metal1 s 754 320 812 329 1 B1
port 3 nsew signal input
rlabel metal1 s 754 292 1364 320 1 B1
port 3 nsew signal input
rlabel metal1 s 754 283 812 292 1 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 1472 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1472 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1472 544
string GDS_END 3645750
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3635170
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 36.800 0.000 
<< end >>
