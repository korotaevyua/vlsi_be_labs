magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1027 203
rect 30 -17 64 21
<< locali >>
rect 371 323 405 493
rect 539 323 573 493
rect 707 323 741 493
rect 875 323 909 493
rect 371 289 909 323
rect 28 215 248 255
rect 858 181 909 289
rect 371 147 909 181
rect 371 51 405 147
rect 539 51 573 147
rect 707 51 741 147
rect 875 51 909 147
<< obsli1 >>
rect 0 527 1104 561
rect 19 323 85 493
rect 119 367 153 527
rect 187 323 253 493
rect 287 367 321 527
rect 439 367 505 527
rect 607 367 673 527
rect 775 367 841 527
rect 19 289 319 323
rect 943 297 1009 527
rect 284 249 319 289
rect 284 215 809 249
rect 284 181 319 215
rect 35 147 319 181
rect 35 51 69 147
rect 103 17 169 113
rect 203 52 237 147
rect 271 17 337 113
rect 439 17 505 113
rect 607 17 673 113
rect 775 17 841 113
rect 943 17 1009 177
rect 0 -17 1104 17
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< labels >>
rlabel locali s 28 215 248 255 6 A
port 1 nsew signal input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 1027 203 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 875 51 909 147 6 X
port 6 nsew signal output
rlabel locali s 707 51 741 147 6 X
port 6 nsew signal output
rlabel locali s 539 51 573 147 6 X
port 6 nsew signal output
rlabel locali s 371 51 405 147 6 X
port 6 nsew signal output
rlabel locali s 371 147 909 181 6 X
port 6 nsew signal output
rlabel locali s 858 181 909 289 6 X
port 6 nsew signal output
rlabel locali s 371 289 909 323 6 X
port 6 nsew signal output
rlabel locali s 875 323 909 493 6 X
port 6 nsew signal output
rlabel locali s 707 323 741 493 6 X
port 6 nsew signal output
rlabel locali s 539 323 573 493 6 X
port 6 nsew signal output
rlabel locali s 371 323 405 493 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3113382
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3104550
<< end >>
