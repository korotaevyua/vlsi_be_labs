magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 827 203
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 177
rect 158 47 188 177
rect 255 47 285 177
rect 372 47 402 177
rect 467 47 497 177
rect 551 47 581 177
rect 635 47 665 177
rect 719 47 749 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 255 297 285 497
rect 371 297 401 497
rect 467 297 497 497
rect 551 297 581 497
rect 635 297 665 497
rect 719 297 749 497
<< ndiff >>
rect 27 101 79 177
rect 27 67 35 101
rect 69 67 79 101
rect 27 47 79 67
rect 109 47 158 177
rect 188 47 255 177
rect 285 47 372 177
rect 402 94 467 177
rect 402 60 421 94
rect 455 60 467 94
rect 402 47 467 60
rect 497 101 551 177
rect 497 67 507 101
rect 541 67 551 101
rect 497 47 551 67
rect 581 94 635 177
rect 581 60 591 94
rect 625 60 635 94
rect 581 47 635 60
rect 665 101 719 177
rect 665 67 675 101
rect 709 67 719 101
rect 665 47 719 67
rect 749 94 801 177
rect 749 60 759 94
rect 793 60 801 94
rect 749 47 801 60
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 297 79 383
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 489 255 497
rect 193 455 207 489
rect 241 455 255 489
rect 193 421 255 455
rect 193 387 207 421
rect 241 387 255 421
rect 193 297 255 387
rect 285 477 371 497
rect 285 443 295 477
rect 329 443 371 477
rect 285 409 371 443
rect 285 375 295 409
rect 329 375 371 409
rect 285 297 371 375
rect 401 489 467 497
rect 401 455 421 489
rect 455 455 467 489
rect 401 421 467 455
rect 401 387 421 421
rect 455 387 467 421
rect 401 297 467 387
rect 497 477 551 497
rect 497 443 507 477
rect 541 443 551 477
rect 497 409 551 443
rect 497 375 507 409
rect 541 375 551 409
rect 497 297 551 375
rect 581 485 635 497
rect 581 451 591 485
rect 625 451 635 485
rect 581 417 635 451
rect 581 383 591 417
rect 625 383 635 417
rect 581 297 635 383
rect 665 477 719 497
rect 665 443 675 477
rect 709 443 719 477
rect 665 409 719 443
rect 665 375 675 409
rect 709 375 719 409
rect 665 297 719 375
rect 749 485 801 497
rect 749 451 759 485
rect 793 451 801 485
rect 749 417 801 451
rect 749 383 759 417
rect 793 383 801 417
rect 749 297 801 383
<< ndiffc >>
rect 35 67 69 101
rect 421 60 455 94
rect 507 67 541 101
rect 591 60 625 94
rect 675 67 709 101
rect 759 60 793 94
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 119 443 153 477
rect 119 375 153 409
rect 207 455 241 489
rect 207 387 241 421
rect 295 443 329 477
rect 295 375 329 409
rect 421 455 455 489
rect 421 387 455 421
rect 507 443 541 477
rect 507 375 541 409
rect 591 451 625 485
rect 591 383 625 417
rect 675 443 709 477
rect 675 375 709 409
rect 759 451 793 485
rect 759 383 793 417
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 255 497 285 523
rect 371 497 401 523
rect 467 497 497 523
rect 551 497 581 523
rect 635 497 665 523
rect 719 497 749 523
rect 79 265 109 297
rect 163 265 193 297
rect 255 265 285 297
rect 371 265 401 297
rect 467 265 497 297
rect 551 265 581 297
rect 635 265 665 297
rect 719 265 749 297
rect 22 249 109 265
rect 22 215 32 249
rect 66 215 109 249
rect 22 199 109 215
rect 79 177 109 199
rect 158 249 212 265
rect 158 215 168 249
rect 202 215 212 249
rect 158 199 212 215
rect 254 249 327 265
rect 254 215 283 249
rect 317 215 327 249
rect 254 199 327 215
rect 371 249 425 265
rect 371 215 381 249
rect 415 215 425 249
rect 158 177 188 199
rect 255 177 285 199
rect 371 193 425 215
rect 467 249 749 265
rect 467 215 531 249
rect 565 215 599 249
rect 633 215 667 249
rect 701 215 749 249
rect 467 199 749 215
rect 372 177 402 193
rect 467 177 497 199
rect 551 177 581 199
rect 635 177 665 199
rect 719 177 749 199
rect 79 21 109 47
rect 158 21 188 47
rect 255 21 285 47
rect 372 21 402 47
rect 467 21 497 47
rect 551 21 581 47
rect 635 21 665 47
rect 719 21 749 47
<< polycont >>
rect 32 215 66 249
rect 168 215 202 249
rect 283 215 317 249
rect 381 215 415 249
rect 531 215 565 249
rect 599 215 633 249
rect 667 215 701 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 21 485 77 527
rect 21 451 35 485
rect 69 451 77 485
rect 21 417 77 451
rect 21 383 35 417
rect 69 383 77 417
rect 21 367 77 383
rect 111 477 153 493
rect 111 443 119 477
rect 111 409 153 443
rect 111 375 119 409
rect 191 489 257 527
rect 191 455 207 489
rect 241 455 257 489
rect 191 421 257 455
rect 191 387 207 421
rect 241 387 257 421
rect 291 477 329 493
rect 291 443 295 477
rect 291 409 329 443
rect 111 333 153 375
rect 291 375 295 409
rect 291 333 329 375
rect 405 489 471 527
rect 405 455 421 489
rect 455 455 471 489
rect 405 421 471 455
rect 405 387 421 421
rect 455 387 471 421
rect 405 371 471 387
rect 507 477 557 493
rect 541 443 557 477
rect 507 409 557 443
rect 541 375 557 409
rect 507 359 557 375
rect 591 485 641 527
rect 625 451 641 485
rect 591 417 641 451
rect 625 383 641 417
rect 591 367 641 383
rect 675 477 709 493
rect 675 409 709 443
rect 743 485 809 527
rect 743 451 759 485
rect 793 451 809 485
rect 743 417 809 451
rect 743 383 759 417
rect 793 383 809 417
rect 25 249 66 331
rect 25 215 32 249
rect 25 153 66 215
rect 100 299 483 333
rect 100 117 134 299
rect 168 249 249 265
rect 202 215 249 249
rect 168 199 249 215
rect 35 101 134 117
rect 69 67 134 101
rect 178 84 249 199
rect 283 249 340 265
rect 317 215 340 249
rect 283 85 340 215
rect 381 249 415 265
rect 449 261 483 299
rect 523 331 557 359
rect 675 349 709 375
rect 675 331 810 349
rect 523 297 810 331
rect 449 249 717 261
rect 449 221 531 249
rect 515 215 531 221
rect 565 215 599 249
rect 633 215 667 249
rect 701 215 717 249
rect 381 187 415 215
rect 381 146 431 187
rect 760 162 810 297
rect 507 128 810 162
rect 405 94 467 110
rect 35 51 134 67
rect 405 60 421 94
rect 455 60 467 94
rect 405 17 467 60
rect 507 101 541 128
rect 675 101 709 128
rect 507 51 541 67
rect 575 60 591 94
rect 625 60 641 94
rect 575 17 641 60
rect 675 51 709 67
rect 743 60 759 94
rect 793 60 809 94
rect 743 17 809 60
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
<< metal1 >>
rect 0 561 828 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 828 561
rect 0 496 828 527
rect 0 17 828 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 828 17
rect 0 -48 828 -17
<< labels >>
flabel locali s 764 153 798 187 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 764 221 798 255 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel locali s 306 85 340 119 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A
port 1 nsew signal input
flabel locali s 214 85 248 119 0 FreeSans 200 0 0 0 B
port 2 nsew signal input
flabel locali s 396 153 430 187 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 764 289 798 323 0 FreeSans 200 0 0 0 X
port 9 nsew signal output
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 and4_4
rlabel metal1 s 0 -48 828 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 828 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 828 544
string GDS_END 3034890
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3027500
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 20.700 0.000 
<< end >>
