magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1602 582
<< pwell >>
rect 834 157 1563 203
rect 1 21 1563 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 351 47 381 131
rect 435 47 465 131
rect 543 47 573 119
rect 629 47 659 119
rect 724 47 754 131
rect 912 47 942 177
rect 1004 47 1034 177
rect 1172 47 1202 177
rect 1360 47 1390 131
rect 1455 47 1485 177
<< scpmoshvt >>
rect 79 363 109 491
rect 163 363 193 491
rect 351 369 381 497
rect 435 369 465 497
rect 531 413 561 497
rect 652 413 682 497
rect 724 413 754 497
rect 912 297 942 497
rect 1004 297 1034 497
rect 1172 297 1202 497
rect 1360 369 1390 497
rect 1455 297 1485 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 119 351 131
rect 299 85 307 119
rect 341 85 351 119
rect 299 47 351 85
rect 381 89 435 131
rect 381 55 391 89
rect 425 55 435 89
rect 381 47 435 55
rect 465 119 515 131
rect 674 119 724 131
rect 465 47 543 119
rect 573 107 629 119
rect 573 73 584 107
rect 618 73 629 107
rect 573 47 629 73
rect 659 47 724 119
rect 754 106 806 131
rect 754 72 764 106
rect 798 72 806 106
rect 754 47 806 72
rect 860 129 912 177
rect 860 95 868 129
rect 902 95 912 129
rect 860 47 912 95
rect 942 47 1004 177
rect 1034 89 1172 177
rect 1034 55 1055 89
rect 1089 55 1125 89
rect 1159 55 1172 89
rect 1034 47 1172 55
rect 1202 119 1254 177
rect 1405 131 1455 177
rect 1202 85 1212 119
rect 1246 85 1254 119
rect 1202 47 1254 85
rect 1308 119 1360 131
rect 1308 85 1316 119
rect 1350 85 1360 119
rect 1308 47 1360 85
rect 1390 93 1455 131
rect 1390 59 1411 93
rect 1445 59 1455 93
rect 1390 47 1455 59
rect 1485 103 1537 177
rect 1485 69 1495 103
rect 1529 69 1537 103
rect 1485 47 1537 69
<< pdiff >>
rect 27 477 79 491
rect 27 443 35 477
rect 69 443 79 477
rect 27 409 79 443
rect 27 375 35 409
rect 69 375 79 409
rect 27 363 79 375
rect 109 461 163 491
rect 109 427 119 461
rect 153 427 163 461
rect 109 363 163 427
rect 193 477 245 491
rect 193 443 203 477
rect 237 443 245 477
rect 193 409 245 443
rect 193 375 203 409
rect 237 375 245 409
rect 193 363 245 375
rect 299 483 351 497
rect 299 449 307 483
rect 341 449 351 483
rect 299 415 351 449
rect 299 381 307 415
rect 341 381 351 415
rect 299 369 351 381
rect 381 485 435 497
rect 381 451 391 485
rect 425 451 435 485
rect 381 417 435 451
rect 381 383 391 417
rect 425 383 435 417
rect 381 369 435 383
rect 465 413 531 497
rect 561 485 652 497
rect 561 451 596 485
rect 630 451 652 485
rect 561 413 652 451
rect 682 413 724 497
rect 754 477 806 497
rect 754 443 764 477
rect 798 443 806 477
rect 754 413 806 443
rect 860 485 912 497
rect 860 451 868 485
rect 902 451 912 485
rect 465 369 515 413
rect 860 297 912 451
rect 942 471 1004 497
rect 942 437 960 471
rect 994 437 1004 471
rect 942 368 1004 437
rect 942 334 960 368
rect 994 334 1004 368
rect 942 297 1004 334
rect 1034 489 1172 497
rect 1034 387 1060 489
rect 1162 387 1172 489
rect 1034 297 1172 387
rect 1202 477 1254 497
rect 1202 443 1212 477
rect 1246 443 1254 477
rect 1202 409 1254 443
rect 1202 375 1212 409
rect 1246 375 1254 409
rect 1202 297 1254 375
rect 1308 450 1360 497
rect 1308 416 1316 450
rect 1350 416 1360 450
rect 1308 369 1360 416
rect 1390 485 1455 497
rect 1390 451 1411 485
rect 1445 451 1455 485
rect 1390 417 1455 451
rect 1390 383 1411 417
rect 1445 383 1455 417
rect 1390 369 1455 383
rect 1405 297 1455 369
rect 1485 477 1537 497
rect 1485 443 1495 477
rect 1529 443 1537 477
rect 1485 409 1537 443
rect 1485 375 1495 409
rect 1529 375 1537 409
rect 1485 297 1537 375
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 307 85 341 119
rect 391 55 425 89
rect 584 73 618 107
rect 764 72 798 106
rect 868 95 902 129
rect 1055 55 1089 89
rect 1125 55 1159 89
rect 1212 85 1246 119
rect 1316 85 1350 119
rect 1411 59 1445 93
rect 1495 69 1529 103
<< pdiffc >>
rect 35 443 69 477
rect 35 375 69 409
rect 119 427 153 461
rect 203 443 237 477
rect 203 375 237 409
rect 307 449 341 483
rect 307 381 341 415
rect 391 451 425 485
rect 391 383 425 417
rect 596 451 630 485
rect 764 443 798 477
rect 868 451 902 485
rect 960 437 994 471
rect 960 334 994 368
rect 1060 387 1162 489
rect 1212 443 1246 477
rect 1212 375 1246 409
rect 1316 416 1350 450
rect 1411 451 1445 485
rect 1411 383 1445 417
rect 1495 443 1529 477
rect 1495 375 1529 409
<< poly >>
rect 79 491 109 517
rect 163 491 193 517
rect 351 497 381 523
rect 435 497 465 523
rect 531 497 561 523
rect 652 497 682 523
rect 724 497 754 523
rect 912 497 942 523
rect 1004 497 1034 523
rect 1172 497 1202 523
rect 1360 497 1390 523
rect 1455 497 1485 523
rect 79 348 109 363
rect 46 318 109 348
rect 46 280 76 318
rect 21 264 76 280
rect 163 274 193 363
rect 21 230 32 264
rect 66 230 76 264
rect 21 214 76 230
rect 118 264 193 274
rect 118 230 134 264
rect 168 230 193 264
rect 351 241 381 369
rect 118 220 193 230
rect 46 176 76 214
rect 46 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 298 225 381 241
rect 298 191 308 225
rect 342 191 381 225
rect 435 219 465 369
rect 531 337 561 413
rect 652 375 682 413
rect 507 321 561 337
rect 603 365 682 375
rect 603 331 619 365
rect 653 331 682 365
rect 603 321 682 331
rect 724 373 754 413
rect 724 357 812 373
rect 724 323 768 357
rect 802 323 812 357
rect 507 287 517 321
rect 551 287 561 321
rect 507 279 561 287
rect 724 307 812 323
rect 507 271 659 279
rect 531 249 659 271
rect 298 175 381 191
rect 351 131 381 175
rect 424 203 478 219
rect 424 169 434 203
rect 468 169 478 203
rect 424 153 478 169
rect 533 191 587 207
rect 533 157 543 191
rect 577 157 587 191
rect 435 131 465 153
rect 533 141 587 157
rect 543 119 573 141
rect 629 119 659 249
rect 724 131 754 307
rect 1360 354 1390 369
rect 1334 324 1390 354
rect 912 265 942 297
rect 1004 265 1034 297
rect 1172 265 1202 297
rect 1334 265 1364 324
rect 1455 265 1485 297
rect 800 249 942 265
rect 800 215 810 249
rect 844 215 942 249
rect 800 199 942 215
rect 984 249 1038 265
rect 984 215 994 249
rect 1028 215 1038 249
rect 984 199 1038 215
rect 1131 249 1364 265
rect 1131 215 1141 249
rect 1175 215 1364 249
rect 1131 199 1364 215
rect 1426 249 1488 265
rect 1426 215 1444 249
rect 1478 215 1488 249
rect 1426 199 1488 215
rect 912 177 942 199
rect 1004 177 1034 199
rect 1172 177 1202 199
rect 1334 176 1364 199
rect 1455 177 1485 199
rect 1334 146 1390 176
rect 1360 131 1390 146
rect 79 21 109 47
rect 163 21 193 47
rect 351 21 381 47
rect 435 21 465 47
rect 543 21 573 47
rect 629 21 659 47
rect 724 21 754 47
rect 912 21 942 47
rect 1004 21 1034 47
rect 1172 21 1202 47
rect 1360 21 1390 47
rect 1455 21 1485 47
<< polycont >>
rect 32 230 66 264
rect 134 230 168 264
rect 308 191 342 225
rect 619 331 653 365
rect 768 323 802 357
rect 517 287 551 321
rect 434 169 468 203
rect 543 157 577 191
rect 810 215 844 249
rect 994 215 1028 249
rect 1141 215 1175 249
rect 1444 215 1478 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 17 477 69 493
rect 17 443 35 477
rect 17 409 69 443
rect 103 461 169 527
rect 103 427 119 461
rect 153 427 169 461
rect 203 477 248 493
rect 391 485 454 527
rect 237 443 248 477
rect 17 375 35 409
rect 203 409 248 443
rect 69 375 156 393
rect 17 359 156 375
rect 17 264 66 325
rect 17 230 32 264
rect 17 197 66 230
rect 122 323 156 359
rect 122 280 156 289
rect 237 391 248 409
rect 203 357 214 375
rect 203 337 248 357
rect 291 449 307 483
rect 341 449 357 483
rect 291 415 357 449
rect 291 381 307 415
rect 341 381 357 415
rect 122 264 168 280
rect 122 230 134 264
rect 122 214 168 230
rect 122 161 156 214
rect 17 127 156 161
rect 17 119 69 127
rect 17 85 35 119
rect 203 119 237 337
rect 291 333 357 381
rect 425 451 454 485
rect 580 451 596 485
rect 630 451 730 485
rect 391 417 454 451
rect 425 383 454 417
rect 391 367 454 383
rect 494 391 551 401
rect 528 357 551 391
rect 291 299 428 333
rect 292 225 358 265
rect 292 191 308 225
rect 342 191 358 225
rect 394 219 428 299
rect 494 321 551 357
rect 494 287 517 321
rect 494 271 551 287
rect 585 365 653 399
rect 585 331 619 365
rect 585 323 653 331
rect 585 289 586 323
rect 620 289 653 323
rect 585 283 653 289
rect 394 203 468 219
rect 585 207 619 283
rect 696 265 730 451
rect 764 477 818 527
rect 798 443 818 477
rect 764 427 818 443
rect 852 485 918 527
rect 1030 489 1178 527
rect 852 451 868 485
rect 902 451 918 485
rect 852 427 918 451
rect 952 471 994 487
rect 952 437 960 471
rect 952 373 994 437
rect 1030 387 1060 489
rect 1162 387 1178 489
rect 1212 477 1276 493
rect 1246 443 1276 477
rect 1212 409 1276 443
rect 768 368 994 373
rect 768 357 960 368
rect 802 334 960 357
rect 1246 375 1276 409
rect 994 334 1175 353
rect 802 323 1175 334
rect 768 307 1175 323
rect 696 249 860 265
rect 696 233 810 249
rect 394 169 434 203
rect 394 157 468 169
rect 17 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 203 69 237 85
rect 307 153 468 157
rect 543 191 619 207
rect 577 157 619 191
rect 307 123 428 153
rect 543 141 619 157
rect 666 215 810 233
rect 844 215 860 249
rect 666 199 860 215
rect 894 249 1091 265
rect 894 215 994 249
rect 1028 215 1091 249
rect 894 199 1091 215
rect 1125 249 1175 307
rect 1125 215 1141 249
rect 307 119 341 123
rect 666 107 700 199
rect 1125 165 1175 215
rect 307 69 341 85
rect 103 17 169 59
rect 375 55 391 89
rect 425 55 441 89
rect 568 73 584 107
rect 618 73 700 107
rect 848 131 1175 165
rect 848 129 908 131
rect 375 17 441 55
rect 748 72 764 106
rect 798 72 814 106
rect 748 17 814 72
rect 848 95 868 129
rect 902 95 908 129
rect 1212 119 1276 375
rect 848 51 908 95
rect 1027 89 1175 97
rect 1027 55 1055 89
rect 1089 55 1125 89
rect 1159 55 1175 89
rect 1027 17 1175 55
rect 1246 85 1276 119
rect 1212 51 1276 85
rect 1316 450 1366 493
rect 1350 416 1366 450
rect 1316 265 1366 416
rect 1402 485 1461 527
rect 1402 451 1411 485
rect 1445 451 1461 485
rect 1402 417 1461 451
rect 1402 383 1411 417
rect 1445 383 1461 417
rect 1402 367 1461 383
rect 1495 477 1547 493
rect 1529 443 1547 477
rect 1495 409 1547 443
rect 1529 375 1547 409
rect 1495 357 1547 375
rect 1316 249 1478 265
rect 1316 215 1444 249
rect 1316 199 1478 215
rect 1316 197 1366 199
rect 1316 119 1350 197
rect 1512 119 1547 357
rect 1495 103 1547 119
rect 1316 51 1350 85
rect 1395 59 1411 93
rect 1445 59 1461 93
rect 1395 17 1461 59
rect 1529 69 1547 103
rect 1495 51 1547 69
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 122 289 156 323
rect 214 375 237 391
rect 237 375 248 391
rect 214 357 248 375
rect 494 357 528 391
rect 586 289 620 323
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
<< metal1 >>
rect 0 561 1564 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1564 561
rect 0 496 1564 527
rect 202 391 260 397
rect 202 357 214 391
rect 248 388 260 391
rect 482 391 540 397
rect 482 388 494 391
rect 248 360 494 388
rect 248 357 260 360
rect 202 351 260 357
rect 482 357 494 360
rect 528 357 540 391
rect 482 351 540 357
rect 110 323 168 329
rect 110 289 122 323
rect 156 320 168 323
rect 574 323 632 329
rect 574 320 586 323
rect 156 292 586 320
rect 156 289 168 292
rect 110 283 168 289
rect 574 289 586 292
rect 620 289 632 323
rect 574 283 632 289
rect 0 17 1564 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1564 17
rect 0 -48 1564 -17
<< labels >>
flabel locali s 958 221 992 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1500 85 1534 119 0 FreeSans 200 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1050 221 1084 255 0 FreeSans 200 0 0 0 RESET_B
port 3 nsew signal input
flabel locali s 1220 289 1254 323 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 310 221 344 255 0 FreeSans 200 0 0 0 D
port 1 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1220 357 1254 391 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 GATE_N
port 2 nsew clock input
flabel locali s 1220 425 1254 459 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1220 85 1254 119 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1500 357 1534 391 0 FreeSans 200 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1220 221 1254 255 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel locali s 1500 425 1534 459 0 FreeSans 200 0 0 0 Q_N
port 9 nsew signal output
flabel locali s 1220 153 1254 187 0 FreeSans 200 0 0 0 Q
port 8 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel metal1 s 47 544 47 544 0 FreeSans 200 0 0 0 VPWR
flabel metal1 s 47 0 47 0 0 FreeSans 200 0 0 0 VGND
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel nwell s 47 544 47 544 0 FreeSans 200 0 0 0 VPB
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
flabel pwell s 47 0 47 0 0 FreeSans 200 0 0 0 VNB
rlabel comment s 0 0 0 0 4 dlrbn_1
rlabel metal1 s 0 -48 1564 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1564 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1564 544
string GDS_END 2683232
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2669476
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
<< end >>
