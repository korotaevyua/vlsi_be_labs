magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 825 157 1103 203
rect 1 21 1103 157
rect 30 -17 64 21
<< locali >>
rect 17 197 66 325
rect 287 191 353 265
rect 1035 334 1087 491
rect 1053 149 1087 334
rect 1035 83 1087 149
<< obsli1 >>
rect 0 527 1104 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 156 393
rect 122 280 156 359
rect 203 337 248 493
rect 122 214 168 280
rect 122 161 156 214
rect 35 127 156 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 237 337
rect 286 333 357 483
rect 391 367 449 527
rect 549 451 721 485
rect 659 421 721 451
rect 755 435 819 527
rect 659 418 724 421
rect 678 417 724 418
rect 678 413 726 417
rect 678 409 729 413
rect 681 407 729 409
rect 686 402 729 407
rect 286 299 423 333
rect 389 247 423 299
rect 489 271 556 401
rect 590 312 657 382
rect 389 157 464 247
rect 590 208 653 312
rect 691 290 729 402
rect 859 373 908 487
rect 763 307 908 373
rect 944 314 1001 527
rect 302 153 464 157
rect 302 123 423 153
rect 512 147 653 208
rect 687 265 729 290
rect 874 265 908 307
rect 687 199 840 265
rect 874 199 1019 265
rect 302 69 341 123
rect 687 107 721 199
rect 874 144 908 199
rect 375 17 441 89
rect 553 73 721 107
rect 755 17 809 109
rect 859 52 908 144
rect 951 17 996 143
rect 0 -17 1104 17
<< metal1 >>
rect 0 496 1104 592
rect 0 -48 1104 48
<< obsm1 >>
rect 202 388 260 397
rect 477 388 535 397
rect 202 360 535 388
rect 202 351 260 360
rect 477 351 535 360
rect 110 320 168 329
rect 578 320 636 329
rect 110 292 636 320
rect 110 283 168 292
rect 578 283 636 292
<< labels >>
rlabel locali s 287 191 353 265 6 D
port 1 nsew signal input
rlabel locali s 17 197 66 325 6 GATE_N
port 2 nsew clock input
rlabel metal1 s 0 -48 1104 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1103 157 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 825 157 1103 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1035 83 1087 149 6 Q
port 7 nsew signal output
rlabel locali s 1053 149 1087 334 6 Q
port 7 nsew signal output
rlabel locali s 1035 334 1087 491 6 Q
port 7 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2844680
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2834078
<< end >>
