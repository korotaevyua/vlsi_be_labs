magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 774 582
<< pwell >>
rect 1 21 735 183
rect 29 -17 63 21
<< obsli1 >>
rect 0 527 736 561
rect 17 309 719 493
rect 17 171 347 275
rect 381 205 719 309
rect 17 17 719 171
rect 0 -17 736 17
<< metal1 >>
rect 0 496 736 592
rect 14 428 722 468
rect 17 416 719 428
rect 0 -48 736 48
<< labels >>
rlabel metal1 s 17 416 719 428 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 14 428 722 468 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -48 736 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 735 183 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 774 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 736 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 736 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2342774
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2338522
<< end >>
