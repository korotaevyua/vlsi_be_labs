magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 590 582
<< pwell >>
rect 157 157 549 203
rect 59 21 549 157
rect 59 17 63 21
rect 29 -17 63 17
<< locali >>
rect 21 195 67 333
rect 209 269 275 491
rect 209 209 316 269
rect 267 159 316 209
rect 352 199 431 269
rect 470 199 528 269
rect 267 53 353 159
rect 389 75 431 199
<< obsli1 >>
rect 0 527 552 561
rect 19 409 71 487
rect 105 445 171 527
rect 19 369 171 409
rect 103 233 171 369
rect 309 345 347 491
rect 381 381 447 527
rect 483 345 517 491
rect 309 305 517 345
rect 103 143 149 233
rect 73 53 149 143
rect 185 17 231 173
rect 465 17 531 163
rect 0 -17 552 17
<< metal1 >>
rect 0 496 552 592
rect 0 -48 552 48
<< labels >>
rlabel locali s 389 75 431 199 6 A1
port 1 nsew signal input
rlabel locali s 352 199 431 269 6 A1
port 1 nsew signal input
rlabel locali s 470 199 528 269 6 A2
port 2 nsew signal input
rlabel locali s 21 195 67 333 6 B1_N
port 3 nsew signal input
rlabel metal1 s 0 -48 552 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 17 8 VNB
port 5 nsew ground bidirectional
rlabel pwell s 59 17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 59 21 549 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 157 157 549 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 590 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 552 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 267 53 353 159 6 Y
port 8 nsew signal output
rlabel locali s 267 159 316 209 6 Y
port 8 nsew signal output
rlabel locali s 209 209 316 269 6 Y
port 8 nsew signal output
rlabel locali s 209 269 275 491 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 552 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3994330
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3988094
<< end >>
