magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 2246 582
<< pwell >>
rect 273 157 457 201
rect 1669 181 2189 203
rect 1386 157 2189 181
rect 1 21 2189 157
rect 29 -17 63 21
<< locali >>
rect 18 195 88 325
rect 354 201 436 325
rect 1785 328 1834 493
rect 1953 328 1987 493
rect 2121 328 2191 493
rect 1785 294 2191 328
rect 2145 177 2191 294
rect 1785 143 2191 177
rect 1785 53 1834 143
rect 1953 53 1987 143
rect 2121 53 2191 143
<< obsli1 >>
rect 0 527 2208 561
rect 35 393 69 493
rect 103 427 169 527
rect 35 359 168 393
rect 122 161 168 359
rect 35 127 168 161
rect 35 69 69 127
rect 103 17 169 93
rect 203 69 248 493
rect 291 427 357 527
rect 391 393 425 493
rect 472 450 638 484
rect 686 451 762 527
rect 286 359 425 393
rect 286 165 320 359
rect 470 315 570 391
rect 286 127 425 165
rect 470 141 514 315
rect 604 281 638 450
rect 798 417 832 475
rect 866 451 932 527
rect 1022 433 1148 483
rect 1184 451 1268 527
rect 1114 417 1148 433
rect 1308 417 1356 475
rect 672 367 942 417
rect 672 315 722 367
rect 824 281 874 313
rect 604 247 874 281
rect 604 239 688 247
rect 550 129 620 203
rect 291 17 357 93
rect 391 61 425 127
rect 654 93 688 239
rect 908 213 942 367
rect 722 147 804 213
rect 862 145 942 213
rect 976 331 1080 393
rect 1114 383 1356 417
rect 1402 389 1468 527
rect 976 179 1010 331
rect 1044 213 1080 295
rect 1114 281 1148 383
rect 1502 353 1536 475
rect 1590 383 1656 485
rect 1502 349 1570 353
rect 1182 315 1570 349
rect 1114 247 1494 281
rect 1164 179 1230 203
rect 976 145 1230 179
rect 485 53 688 93
rect 722 17 804 105
rect 862 59 912 145
rect 948 17 1016 109
rect 1264 95 1298 247
rect 1428 235 1494 247
rect 1332 201 1398 213
rect 1332 147 1464 201
rect 1528 136 1570 315
rect 1128 61 1298 95
rect 1334 17 1466 113
rect 1502 70 1570 136
rect 1606 255 1656 383
rect 1692 367 1749 527
rect 1868 362 1919 527
rect 2021 362 2087 527
rect 1606 211 2111 255
rect 1606 69 1656 211
rect 1692 17 1749 109
rect 1868 17 1919 109
rect 2021 17 2087 109
rect 0 -17 2208 17
<< metal1 >>
rect 0 496 2208 592
rect 753 184 811 193
rect 1397 184 1455 193
rect 753 156 1455 184
rect 753 147 811 156
rect 1397 147 1455 156
rect 0 -48 2208 48
<< obsm1 >>
rect 111 388 169 397
rect 477 388 535 397
rect 1029 388 1087 397
rect 111 360 1087 388
rect 111 351 169 360
rect 477 351 535 360
rect 1029 351 1087 360
rect 1033 252 1091 261
rect 584 224 1091 252
rect 584 193 627 224
rect 1033 215 1091 224
rect 201 184 259 193
rect 569 184 627 193
rect 201 156 627 184
rect 201 147 259 156
rect 569 147 627 156
<< labels >>
rlabel locali s 18 195 88 325 6 CLK
port 1 nsew clock input
rlabel locali s 354 201 436 325 6 D
port 2 nsew signal input
rlabel metal1 s 1397 147 1455 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 147 811 156 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 156 1455 184 6 SET_B
port 3 nsew signal input
rlabel metal1 s 1397 184 1455 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 753 184 811 193 6 SET_B
port 3 nsew signal input
rlabel metal1 s 0 -48 2208 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 2189 157 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1386 157 2189 181 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1669 181 2189 203 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 273 157 457 201 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 2246 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 2208 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 2121 53 2191 143 6 Q
port 8 nsew signal output
rlabel locali s 1953 53 1987 143 6 Q
port 8 nsew signal output
rlabel locali s 1785 53 1834 143 6 Q
port 8 nsew signal output
rlabel locali s 1785 143 2191 177 6 Q
port 8 nsew signal output
rlabel locali s 2145 177 2191 294 6 Q
port 8 nsew signal output
rlabel locali s 1785 294 2191 328 6 Q
port 8 nsew signal output
rlabel locali s 2121 328 2191 493 6 Q
port 8 nsew signal output
rlabel locali s 1953 328 1987 493 6 Q
port 8 nsew signal output
rlabel locali s 1785 328 1834 493 6 Q
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 2208 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2564738
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2547064
<< end >>
