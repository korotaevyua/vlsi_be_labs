magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1142 582
<< pwell >>
rect 1 21 1103 183
rect 29 -17 63 21
<< obsli1 >>
rect 0 527 1104 561
rect 17 309 1086 493
rect 17 171 533 275
rect 567 205 1086 309
rect 17 17 1086 171
rect 0 -17 1104 17
<< metal1 >>
rect 0 496 1104 592
rect 14 428 1090 468
rect 17 416 1087 428
rect 0 -48 1104 48
<< labels >>
rlabel metal1 s 17 416 1087 428 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 14 428 1090 468 6 KAPWR
port 1 nsew power bidirectional abutment
rlabel metal1 s 0 -48 1104 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 3 nsew ground bidirectional
rlabel pwell s 1 21 1103 183 6 VNB
port 3 nsew ground bidirectional
rlabel nwell s -38 261 1142 582 6 VPB
port 4 nsew power bidirectional
rlabel metal1 s 0 496 1104 592 6 VPWR
port 5 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1104 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2338454
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2333338
<< end >>
