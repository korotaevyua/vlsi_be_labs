magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 406 582
<< pwell >>
rect 6 21 366 157
rect 29 -17 63 21
<< locali >>
rect 193 336 260 493
rect 17 191 83 323
rect 121 268 155 329
rect 193 302 269 336
rect 121 220 201 268
rect 235 225 269 302
rect 303 271 346 337
rect 235 191 348 225
rect 291 56 348 191
<< obsli1 >>
rect 0 527 368 561
rect 29 365 95 527
rect 294 371 345 527
rect 24 123 257 157
rect 24 56 76 123
rect 110 17 176 89
rect 210 56 257 123
rect 0 -17 368 17
<< metal1 >>
rect 0 496 368 592
rect 0 -48 368 48
<< labels >>
rlabel locali s 17 191 83 323 6 A1
port 1 nsew signal input
rlabel locali s 121 220 201 268 6 A2
port 2 nsew signal input
rlabel locali s 121 268 155 329 6 A2
port 2 nsew signal input
rlabel locali s 303 271 346 337 6 B1
port 3 nsew signal input
rlabel metal1 s 0 -48 368 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 29 -17 63 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 6 21 366 157 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 406 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 368 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 291 56 348 191 6 Y
port 8 nsew signal output
rlabel locali s 235 191 348 225 6 Y
port 8 nsew signal output
rlabel locali s 235 225 269 302 6 Y
port 8 nsew signal output
rlabel locali s 193 302 269 336 6 Y
port 8 nsew signal output
rlabel locali s 193 336 260 493 6 Y
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 368 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1286826
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1282564
<< end >>
