magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1878 582
<< pwell >>
rect 1 21 1839 203
rect 30 -17 64 21
<< locali >>
rect 103 267 169 483
rect 271 313 337 483
rect 271 267 310 313
rect 103 213 310 267
rect 103 63 169 213
rect 271 165 310 213
rect 271 63 337 165
rect 842 301 1362 335
rect 842 249 876 301
rect 664 215 876 249
rect 910 233 944 265
rect 910 199 1091 233
rect 1125 199 1159 301
rect 1316 265 1362 301
rect 1057 175 1091 199
rect 1057 169 1099 175
rect 1057 165 1107 169
rect 1217 165 1263 265
rect 1316 199 1411 265
rect 1519 317 1553 483
rect 1681 317 1737 483
rect 1519 283 1737 317
rect 1057 146 1263 165
rect 1681 181 1737 283
rect 1059 144 1263 146
rect 1062 142 1263 144
rect 1064 139 1263 142
rect 1067 135 1263 139
rect 1069 131 1263 135
rect 1519 147 1737 181
rect 1519 63 1569 147
rect 1681 63 1737 147
<< obsli1 >>
rect 0 527 1840 561
rect 27 299 69 527
rect 203 303 237 527
rect 371 299 473 527
rect 554 387 588 471
rect 638 421 672 527
rect 706 441 866 475
rect 1048 441 1114 527
rect 706 387 740 441
rect 1167 405 1201 471
rect 1235 441 1301 527
rect 1335 405 1369 471
rect 1411 441 1477 527
rect 516 353 740 387
rect 774 371 1479 405
rect 516 249 550 353
rect 774 319 808 371
rect 344 215 550 249
rect 27 17 69 177
rect 203 17 237 177
rect 371 17 419 177
rect 516 163 550 215
rect 584 285 808 319
rect 584 199 618 285
rect 1445 249 1479 371
rect 1587 351 1645 527
rect 1771 299 1813 527
rect 1445 215 1645 249
rect 516 129 609 163
rect 643 129 1023 163
rect 1445 163 1479 215
rect 643 95 677 129
rect 454 61 677 95
rect 711 17 782 93
rect 816 69 850 129
rect 984 117 1023 129
rect 1341 129 1479 163
rect 884 17 950 93
rect 984 51 1038 117
rect 1341 93 1375 129
rect 1077 17 1143 93
rect 1235 59 1375 93
rect 1411 17 1477 93
rect 1603 17 1645 113
rect 1771 17 1813 177
rect 0 -17 1840 17
<< metal1 >>
rect 0 496 1840 592
rect 0 -48 1840 48
<< labels >>
rlabel locali s 1316 199 1411 265 6 A
port 1 nsew signal input
rlabel locali s 1316 265 1362 301 6 A
port 1 nsew signal input
rlabel locali s 1125 199 1159 301 6 A
port 1 nsew signal input
rlabel locali s 664 215 876 249 6 A
port 1 nsew signal input
rlabel locali s 842 249 876 301 6 A
port 1 nsew signal input
rlabel locali s 842 301 1362 335 6 A
port 1 nsew signal input
rlabel locali s 1069 131 1263 135 6 B
port 2 nsew signal input
rlabel locali s 1067 135 1263 139 6 B
port 2 nsew signal input
rlabel locali s 1064 139 1263 142 6 B
port 2 nsew signal input
rlabel locali s 1062 142 1263 144 6 B
port 2 nsew signal input
rlabel locali s 1059 144 1263 146 6 B
port 2 nsew signal input
rlabel locali s 1057 146 1263 165 6 B
port 2 nsew signal input
rlabel locali s 1217 165 1263 265 6 B
port 2 nsew signal input
rlabel locali s 1057 165 1107 169 6 B
port 2 nsew signal input
rlabel locali s 1057 169 1099 175 6 B
port 2 nsew signal input
rlabel locali s 1057 175 1091 199 6 B
port 2 nsew signal input
rlabel locali s 910 199 1091 233 6 B
port 2 nsew signal input
rlabel locali s 910 233 944 265 6 B
port 2 nsew signal input
rlabel metal1 s 0 -48 1840 48 8 VGND
port 3 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 4 nsew ground bidirectional
rlabel pwell s 1 21 1839 203 6 VNB
port 4 nsew ground bidirectional
rlabel nwell s -38 261 1878 582 6 VPB
port 5 nsew power bidirectional
rlabel metal1 s 0 496 1840 592 6 VPWR
port 6 nsew power bidirectional abutment
rlabel locali s 1681 63 1737 147 6 COUT
port 7 nsew signal output
rlabel locali s 1519 63 1569 147 6 COUT
port 7 nsew signal output
rlabel locali s 1519 147 1737 181 6 COUT
port 7 nsew signal output
rlabel locali s 1681 181 1737 283 6 COUT
port 7 nsew signal output
rlabel locali s 1519 283 1737 317 6 COUT
port 7 nsew signal output
rlabel locali s 1681 317 1737 483 6 COUT
port 7 nsew signal output
rlabel locali s 1519 317 1553 483 6 COUT
port 7 nsew signal output
rlabel locali s 271 63 337 165 6 SUM
port 8 nsew signal output
rlabel locali s 271 165 310 213 6 SUM
port 8 nsew signal output
rlabel locali s 103 63 169 213 6 SUM
port 8 nsew signal output
rlabel locali s 103 213 310 267 6 SUM
port 8 nsew signal output
rlabel locali s 271 267 310 313 6 SUM
port 8 nsew signal output
rlabel locali s 271 313 337 483 6 SUM
port 8 nsew signal output
rlabel locali s 103 267 169 483 6 SUM
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1840 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 2190846
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 2176828
<< end >>
