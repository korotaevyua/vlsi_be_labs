magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 958 582
<< pwell >>
rect 98 157 366 203
rect 1 21 919 157
rect 30 -17 64 21
<< locali >>
rect 30 199 66 327
rect 198 309 264 343
rect 203 51 248 309
rect 582 84 635 255
rect 670 85 731 281
rect 765 153 835 261
<< obsli1 >>
rect 0 527 920 561
rect 35 411 69 493
rect 103 451 169 527
rect 298 451 432 527
rect 479 417 513 493
rect 547 451 615 527
rect 649 417 683 493
rect 751 451 817 527
rect 851 417 903 493
rect 35 377 385 411
rect 100 161 134 377
rect 35 127 134 161
rect 35 51 69 127
rect 103 17 169 93
rect 351 265 385 377
rect 447 383 683 417
rect 717 383 903 417
rect 283 161 317 265
rect 351 199 413 265
rect 447 161 481 383
rect 717 349 751 383
rect 515 315 751 349
rect 515 280 549 315
rect 283 127 481 161
rect 282 17 348 93
rect 402 51 436 127
rect 869 117 903 383
rect 767 17 817 117
rect 851 51 903 117
rect 0 -17 920 17
<< metal1 >>
rect 0 496 920 592
rect 0 -48 920 48
<< labels >>
rlabel locali s 30 199 66 327 6 A_N
port 1 nsew signal input
rlabel locali s 765 153 835 261 6 B_N
port 2 nsew signal input
rlabel locali s 582 84 635 255 6 C
port 3 nsew signal input
rlabel locali s 670 85 731 281 6 D
port 4 nsew signal input
rlabel metal1 s 0 -48 920 48 8 VGND
port 5 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 1 21 919 157 6 VNB
port 6 nsew ground bidirectional
rlabel pwell s 98 157 366 203 6 VNB
port 6 nsew ground bidirectional
rlabel nwell s -38 261 958 582 6 VPB
port 7 nsew power bidirectional
rlabel metal1 s 0 496 920 592 6 VPWR
port 8 nsew power bidirectional abutment
rlabel locali s 203 51 248 309 6 X
port 9 nsew signal output
rlabel locali s 198 309 264 343 6 X
port 9 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 920 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 3074894
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3066958
<< end >>
