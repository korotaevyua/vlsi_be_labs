magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 35 21 643 203
rect 35 17 64 21
rect 30 -17 64 17
<< scnmos >>
rect 114 47 144 177
rect 200 47 230 177
rect 298 47 328 177
rect 428 47 458 177
rect 534 47 564 177
<< scpmoshvt >>
rect 80 297 110 497
rect 166 297 196 497
rect 356 297 386 497
rect 442 297 472 497
rect 535 297 565 497
<< ndiff >>
rect 61 93 114 177
rect 61 59 69 93
rect 103 59 114 93
rect 61 47 114 59
rect 144 101 200 177
rect 144 67 155 101
rect 189 67 200 101
rect 144 47 200 67
rect 230 89 298 177
rect 230 55 241 89
rect 275 55 298 89
rect 230 47 298 55
rect 328 101 428 177
rect 328 67 339 101
rect 373 67 428 101
rect 328 47 428 67
rect 458 47 534 177
rect 564 93 617 177
rect 564 59 575 93
rect 609 59 617 93
rect 564 47 617 59
<< pdiff >>
rect 27 485 80 497
rect 27 451 35 485
rect 69 451 80 485
rect 27 386 80 451
rect 27 352 35 386
rect 69 352 80 386
rect 27 297 80 352
rect 110 477 166 497
rect 110 443 121 477
rect 155 443 166 477
rect 110 382 166 443
rect 110 348 121 382
rect 155 348 166 382
rect 110 297 166 348
rect 196 485 249 497
rect 196 451 207 485
rect 241 451 249 485
rect 196 297 249 451
rect 303 477 356 497
rect 303 443 311 477
rect 345 443 356 477
rect 303 393 356 443
rect 303 359 311 393
rect 345 359 356 393
rect 303 297 356 359
rect 386 477 442 497
rect 386 443 397 477
rect 431 443 442 477
rect 386 387 442 443
rect 386 353 397 387
rect 431 353 442 387
rect 386 297 442 353
rect 472 485 535 497
rect 472 451 487 485
rect 521 451 535 485
rect 472 297 535 451
rect 565 477 617 497
rect 565 443 575 477
rect 609 443 617 477
rect 565 387 617 443
rect 565 353 575 387
rect 609 353 617 387
rect 565 297 617 353
<< ndiffc >>
rect 69 59 103 93
rect 155 67 189 101
rect 241 55 275 89
rect 339 67 373 101
rect 575 59 609 93
<< pdiffc >>
rect 35 451 69 485
rect 35 352 69 386
rect 121 443 155 477
rect 121 348 155 382
rect 207 451 241 485
rect 311 443 345 477
rect 311 359 345 393
rect 397 443 431 477
rect 397 353 431 387
rect 487 451 521 485
rect 575 443 609 477
rect 575 353 609 387
<< poly >>
rect 80 497 110 523
rect 166 497 196 523
rect 356 497 386 523
rect 442 497 472 523
rect 535 497 565 523
rect 80 229 110 297
rect 166 265 196 297
rect 356 265 386 297
rect 442 265 472 297
rect 166 249 250 265
rect 166 229 200 249
rect 80 215 200 229
rect 234 215 250 249
rect 80 199 250 215
rect 298 249 386 265
rect 298 215 314 249
rect 348 215 386 249
rect 298 199 386 215
rect 428 249 492 265
rect 428 215 448 249
rect 482 215 492 249
rect 535 261 565 297
rect 535 249 612 261
rect 535 227 562 249
rect 428 199 492 215
rect 534 215 562 227
rect 596 215 612 249
rect 534 203 612 215
rect 534 201 566 203
rect 114 177 144 199
rect 200 177 230 199
rect 298 177 328 199
rect 428 177 458 199
rect 534 177 564 201
rect 114 21 144 47
rect 200 21 230 47
rect 298 21 328 47
rect 428 21 458 47
rect 534 21 564 47
<< polycont >>
rect 200 215 234 249
rect 314 215 348 249
rect 448 215 482 249
rect 562 215 596 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 19 485 77 527
rect 19 451 35 485
rect 69 451 77 485
rect 19 386 77 451
rect 19 352 35 386
rect 69 352 77 386
rect 19 333 77 352
rect 111 477 157 493
rect 111 443 121 477
rect 155 443 157 477
rect 191 485 257 527
rect 191 451 207 485
rect 241 451 257 485
rect 191 444 257 451
rect 295 477 358 493
rect 111 382 157 443
rect 295 443 311 477
rect 345 443 358 477
rect 295 393 358 443
rect 295 384 311 393
rect 111 348 121 382
rect 155 348 157 382
rect 111 165 157 348
rect 191 359 311 384
rect 345 359 358 393
rect 191 338 358 359
rect 392 477 437 493
rect 392 443 397 477
rect 431 443 437 477
rect 392 387 437 443
rect 471 485 537 527
rect 471 451 487 485
rect 521 451 537 485
rect 471 425 537 451
rect 571 477 615 493
rect 571 443 575 477
rect 609 443 615 477
rect 571 387 615 443
rect 392 353 397 387
rect 431 353 575 387
rect 609 353 615 387
rect 191 249 259 338
rect 392 334 615 353
rect 191 215 200 249
rect 234 215 259 249
rect 191 199 259 215
rect 293 249 358 282
rect 293 215 314 249
rect 348 215 358 249
rect 293 199 358 215
rect 448 249 524 265
rect 482 215 524 249
rect 225 165 259 199
rect 111 127 191 165
rect 225 131 373 165
rect 153 101 191 127
rect 53 59 69 93
rect 103 59 119 93
rect 53 17 119 59
rect 153 67 155 101
rect 189 67 191 101
rect 335 101 373 131
rect 153 51 191 67
rect 225 55 241 89
rect 275 55 291 89
rect 225 17 291 55
rect 335 67 339 101
rect 448 73 524 215
rect 562 249 625 265
rect 596 215 625 249
rect 562 150 625 215
rect 561 93 627 113
rect 335 51 373 67
rect 561 59 575 93
rect 609 59 627 93
rect 561 17 627 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 122 425 156 459 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel locali s 306 221 340 255 0 FreeSans 340 0 0 0 B1
port 3 nsew signal input
flabel locali s 490 153 524 187 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 582 221 616 255 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 490 85 524 119 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a21o_2
rlabel metal1 s 0 -48 644 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 4022166
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 4016612
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
