magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1694 582
<< pwell >>
rect 506 157 715 203
rect 1019 157 1646 203
rect 1 21 1646 157
rect 30 -17 64 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 260 47 290 119
rect 365 47 395 119
rect 487 47 517 131
rect 607 47 637 177
rect 795 47 825 131
rect 879 47 909 131
rect 1097 47 1127 177
rect 1169 47 1199 177
rect 1276 47 1306 177
rect 1360 47 1390 177
rect 1444 47 1474 177
rect 1528 47 1558 177
<< scpmoshvt >>
rect 79 369 109 497
rect 151 369 181 497
rect 257 413 287 497
rect 353 413 383 497
rect 471 413 501 497
rect 607 297 637 497
rect 795 303 825 431
rect 905 303 935 431
rect 1097 297 1127 497
rect 1181 297 1211 497
rect 1276 297 1306 497
rect 1360 297 1390 497
rect 1444 297 1474 497
rect 1528 297 1558 497
<< ndiff >>
rect 27 103 79 131
rect 27 69 35 103
rect 69 69 79 103
rect 27 47 79 69
rect 109 89 163 131
rect 109 55 119 89
rect 153 55 163 89
rect 109 47 163 55
rect 193 119 245 131
rect 532 131 607 177
rect 437 119 487 131
rect 193 101 260 119
rect 193 67 203 101
rect 237 67 260 101
rect 193 47 260 67
rect 290 89 365 119
rect 290 55 310 89
rect 344 55 365 89
rect 290 47 365 55
rect 395 47 487 119
rect 517 119 607 131
rect 517 85 546 119
rect 580 85 607 119
rect 517 47 607 85
rect 637 101 689 177
rect 637 67 647 101
rect 681 67 689 101
rect 637 47 689 67
rect 743 110 795 131
rect 743 76 751 110
rect 785 76 795 110
rect 743 47 795 76
rect 825 89 879 131
rect 825 55 835 89
rect 869 55 879 89
rect 825 47 879 55
rect 909 110 961 131
rect 909 76 919 110
rect 953 76 961 110
rect 909 47 961 76
rect 1045 109 1097 177
rect 1045 75 1053 109
rect 1087 75 1097 109
rect 1045 47 1097 75
rect 1127 47 1169 177
rect 1199 89 1276 177
rect 1199 55 1216 89
rect 1250 55 1276 89
rect 1199 47 1276 55
rect 1306 89 1360 177
rect 1306 55 1316 89
rect 1350 55 1360 89
rect 1306 47 1360 55
rect 1390 93 1444 177
rect 1390 59 1400 93
rect 1434 59 1444 93
rect 1390 47 1444 59
rect 1474 101 1528 177
rect 1474 67 1484 101
rect 1518 67 1528 101
rect 1474 47 1528 67
rect 1558 161 1620 177
rect 1558 127 1578 161
rect 1612 127 1620 161
rect 1558 93 1620 127
rect 1558 59 1578 93
rect 1612 59 1620 93
rect 1558 47 1620 59
<< pdiff >>
rect 27 485 79 497
rect 27 451 35 485
rect 69 451 79 485
rect 27 417 79 451
rect 27 383 35 417
rect 69 383 79 417
rect 27 369 79 383
rect 109 369 151 497
rect 181 475 257 497
rect 181 441 202 475
rect 236 441 257 475
rect 181 413 257 441
rect 287 480 353 497
rect 287 446 303 480
rect 337 446 353 480
rect 287 413 353 446
rect 383 413 471 497
rect 501 489 607 497
rect 501 455 542 489
rect 576 455 607 489
rect 501 413 607 455
rect 181 369 242 413
rect 557 297 607 413
rect 637 458 689 497
rect 637 424 647 458
rect 681 424 689 458
rect 840 485 890 497
rect 840 451 848 485
rect 882 451 890 485
rect 840 431 890 451
rect 1041 489 1097 497
rect 1041 455 1053 489
rect 1087 455 1097 489
rect 637 297 689 424
rect 743 349 795 431
rect 743 315 751 349
rect 785 315 795 349
rect 743 303 795 315
rect 825 303 905 431
rect 935 349 987 431
rect 935 315 945 349
rect 979 315 987 349
rect 935 303 987 315
rect 1041 297 1097 455
rect 1127 442 1181 497
rect 1127 408 1137 442
rect 1171 408 1181 442
rect 1127 297 1181 408
rect 1211 489 1276 497
rect 1211 455 1227 489
rect 1261 455 1276 489
rect 1211 297 1276 455
rect 1306 448 1360 497
rect 1306 414 1316 448
rect 1350 414 1360 448
rect 1306 380 1360 414
rect 1306 346 1316 380
rect 1350 346 1360 380
rect 1306 297 1360 346
rect 1390 485 1444 497
rect 1390 451 1400 485
rect 1434 451 1444 485
rect 1390 417 1444 451
rect 1390 383 1400 417
rect 1434 383 1444 417
rect 1390 297 1444 383
rect 1474 448 1528 497
rect 1474 414 1484 448
rect 1518 414 1528 448
rect 1474 380 1528 414
rect 1474 346 1484 380
rect 1518 346 1528 380
rect 1474 297 1528 346
rect 1558 485 1620 497
rect 1558 451 1578 485
rect 1612 451 1620 485
rect 1558 417 1620 451
rect 1558 383 1578 417
rect 1612 383 1620 417
rect 1558 349 1620 383
rect 1558 315 1578 349
rect 1612 315 1620 349
rect 1558 297 1620 315
<< ndiffc >>
rect 35 69 69 103
rect 119 55 153 89
rect 203 67 237 101
rect 310 55 344 89
rect 546 85 580 119
rect 647 67 681 101
rect 751 76 785 110
rect 835 55 869 89
rect 919 76 953 110
rect 1053 75 1087 109
rect 1216 55 1250 89
rect 1316 55 1350 89
rect 1400 59 1434 93
rect 1484 67 1518 101
rect 1578 127 1612 161
rect 1578 59 1612 93
<< pdiffc >>
rect 35 451 69 485
rect 35 383 69 417
rect 202 441 236 475
rect 303 446 337 480
rect 542 455 576 489
rect 647 424 681 458
rect 848 451 882 485
rect 1053 455 1087 489
rect 751 315 785 349
rect 945 315 979 349
rect 1137 408 1171 442
rect 1227 455 1261 489
rect 1316 414 1350 448
rect 1316 346 1350 380
rect 1400 451 1434 485
rect 1400 383 1434 417
rect 1484 414 1518 448
rect 1484 346 1518 380
rect 1578 451 1612 485
rect 1578 383 1612 417
rect 1578 315 1612 349
<< poly >>
rect 79 497 109 523
rect 151 497 181 523
rect 257 497 287 523
rect 353 497 383 523
rect 471 497 501 523
rect 607 497 637 523
rect 79 265 109 369
rect 22 249 109 265
rect 22 215 32 249
rect 66 215 109 249
rect 22 199 109 215
rect 151 265 181 369
rect 257 273 287 413
rect 353 381 383 413
rect 471 381 501 413
rect 329 365 383 381
rect 329 331 339 365
rect 373 331 383 365
rect 329 315 383 331
rect 465 365 519 381
rect 465 331 475 365
rect 509 331 519 365
rect 465 315 519 331
rect 151 249 215 265
rect 151 215 171 249
rect 205 215 215 249
rect 257 243 395 273
rect 151 199 215 215
rect 365 207 395 243
rect 79 131 109 199
rect 163 131 193 199
rect 257 191 323 201
rect 257 157 273 191
rect 307 157 323 191
rect 257 147 323 157
rect 365 191 419 207
rect 365 157 375 191
rect 409 157 419 191
rect 260 119 290 147
rect 365 141 419 157
rect 365 119 395 141
rect 487 131 517 315
rect 795 431 825 523
rect 905 431 935 523
rect 1097 497 1127 523
rect 1181 497 1211 523
rect 1276 497 1306 523
rect 1360 497 1390 523
rect 1444 497 1474 523
rect 1528 497 1558 523
rect 607 265 637 297
rect 795 265 825 303
rect 905 265 935 303
rect 1097 265 1127 297
rect 1181 265 1211 297
rect 559 249 637 265
rect 559 215 569 249
rect 603 215 637 249
rect 559 199 637 215
rect 787 255 853 265
rect 787 221 803 255
rect 837 221 853 255
rect 787 211 853 221
rect 905 249 989 265
rect 905 215 945 249
rect 979 215 989 249
rect 607 177 637 199
rect 795 131 825 211
rect 905 176 989 215
rect 1051 249 1127 265
rect 1051 215 1061 249
rect 1095 215 1127 249
rect 1051 199 1127 215
rect 1097 177 1127 199
rect 1169 249 1223 265
rect 1169 215 1179 249
rect 1213 215 1223 249
rect 1169 199 1223 215
rect 1276 259 1306 297
rect 1360 259 1390 297
rect 1444 259 1474 297
rect 1528 259 1558 297
rect 1276 249 1558 259
rect 1276 215 1292 249
rect 1326 215 1558 249
rect 1276 205 1558 215
rect 1169 177 1199 199
rect 1276 177 1306 205
rect 1360 177 1390 205
rect 1444 177 1474 205
rect 1528 177 1558 205
rect 879 146 989 176
rect 879 131 909 146
rect 79 21 109 47
rect 163 21 193 47
rect 260 21 290 47
rect 365 21 395 47
rect 487 21 517 47
rect 607 21 637 47
rect 795 21 825 47
rect 879 21 909 47
rect 1097 21 1127 47
rect 1169 21 1199 47
rect 1276 21 1306 47
rect 1360 21 1390 47
rect 1444 21 1474 47
rect 1528 21 1558 47
<< polycont >>
rect 32 215 66 249
rect 339 331 373 365
rect 475 331 509 365
rect 171 215 205 249
rect 273 157 307 191
rect 375 157 409 191
rect 569 215 603 249
rect 803 221 837 255
rect 945 215 979 249
rect 1061 215 1095 249
rect 1179 215 1213 249
rect 1292 215 1326 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 17 485 69 527
rect 17 451 35 485
rect 17 417 69 451
rect 17 383 35 417
rect 17 367 69 383
rect 103 475 252 493
rect 103 441 202 475
rect 236 441 252 475
rect 103 425 252 441
rect 286 480 441 493
rect 286 446 303 480
rect 337 446 441 480
rect 286 425 441 446
rect 17 249 69 333
rect 17 215 32 249
rect 66 215 69 249
rect 17 191 69 215
rect 103 157 137 425
rect 171 289 248 391
rect 282 365 373 391
rect 282 331 339 365
rect 282 323 373 331
rect 282 289 306 323
rect 340 289 373 323
rect 171 249 239 289
rect 282 265 373 289
rect 205 215 239 249
rect 171 191 239 215
rect 273 241 373 265
rect 407 275 441 425
rect 475 489 603 527
rect 475 455 542 489
rect 576 455 603 489
rect 475 415 603 455
rect 637 458 681 493
rect 637 424 647 458
rect 719 489 1103 527
rect 719 485 1053 489
rect 719 451 848 485
rect 882 455 1053 485
rect 1087 455 1103 489
rect 882 451 1103 455
rect 637 417 681 424
rect 1137 442 1171 493
rect 1211 489 1277 527
rect 1211 455 1227 489
rect 1261 455 1277 489
rect 1211 451 1277 455
rect 637 383 1103 417
rect 637 381 681 383
rect 475 365 681 381
rect 509 331 681 365
rect 475 327 681 331
rect 475 315 509 327
rect 407 249 603 275
rect 407 241 569 249
rect 273 191 341 241
rect 466 215 569 241
rect 307 157 341 191
rect 17 123 239 157
rect 273 141 341 157
rect 375 191 432 207
rect 409 187 432 191
rect 375 153 398 157
rect 375 141 432 153
rect 466 199 603 215
rect 17 103 69 123
rect 17 69 35 103
rect 203 101 239 123
rect 466 107 500 199
rect 17 51 69 69
rect 103 55 119 89
rect 153 55 169 89
rect 103 17 169 55
rect 237 67 239 101
rect 203 51 239 67
rect 273 89 500 107
rect 273 55 310 89
rect 344 55 500 89
rect 273 51 500 55
rect 534 119 603 165
rect 534 85 546 119
rect 580 85 603 119
rect 534 17 603 85
rect 637 101 681 327
rect 637 67 647 101
rect 637 51 681 67
rect 719 315 751 349
rect 785 315 801 349
rect 835 323 945 349
rect 719 187 753 315
rect 835 289 862 323
rect 896 315 945 323
rect 979 315 995 349
rect 896 299 995 315
rect 835 255 896 289
rect 787 221 803 255
rect 837 221 896 255
rect 719 153 770 187
rect 838 157 896 221
rect 945 255 989 265
rect 945 249 954 255
rect 988 221 989 255
rect 979 215 989 221
rect 945 199 989 215
rect 1033 249 1103 383
rect 1316 448 1366 493
rect 1171 408 1282 417
rect 1137 299 1282 408
rect 1033 215 1061 249
rect 1095 215 1103 249
rect 1033 199 1103 215
rect 1137 255 1213 265
rect 1137 221 1142 255
rect 1176 249 1213 255
rect 1176 221 1179 249
rect 1137 215 1179 221
rect 1137 199 1213 215
rect 1248 263 1282 299
rect 1350 414 1366 448
rect 1316 380 1366 414
rect 1350 346 1366 380
rect 1400 485 1450 527
rect 1434 451 1450 485
rect 1400 417 1450 451
rect 1434 383 1450 417
rect 1400 365 1450 383
rect 1484 448 1544 493
rect 1518 414 1544 448
rect 1484 380 1544 414
rect 1316 331 1366 346
rect 1518 346 1544 380
rect 1316 297 1444 331
rect 1410 263 1444 297
rect 1484 263 1544 346
rect 1578 485 1639 527
rect 1612 451 1639 485
rect 1578 417 1639 451
rect 1612 383 1639 417
rect 1578 349 1639 383
rect 1612 315 1639 349
rect 1578 297 1639 315
rect 1248 249 1376 263
rect 1248 215 1292 249
rect 1326 215 1376 249
rect 1248 211 1376 215
rect 1410 211 1639 263
rect 1248 157 1282 211
rect 1410 177 1444 211
rect 719 110 785 153
rect 838 123 969 157
rect 719 76 751 110
rect 919 110 969 123
rect 719 51 785 76
rect 819 55 835 89
rect 869 55 885 89
rect 819 17 885 55
rect 953 76 969 110
rect 919 51 969 76
rect 1003 123 1282 157
rect 1316 143 1444 177
rect 1003 109 1087 123
rect 1003 75 1053 109
rect 1316 89 1366 143
rect 1003 51 1087 75
rect 1121 55 1216 89
rect 1250 55 1266 89
rect 1121 17 1266 55
rect 1300 55 1316 89
rect 1350 55 1366 89
rect 1300 51 1366 55
rect 1400 93 1450 109
rect 1434 59 1450 93
rect 1400 17 1450 59
rect 1484 101 1544 211
rect 1518 67 1544 101
rect 1484 51 1544 67
rect 1578 161 1639 177
rect 1612 127 1639 161
rect 1578 93 1639 127
rect 1612 59 1639 93
rect 1578 17 1639 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 306 289 340 323
rect 398 157 409 187
rect 409 157 432 187
rect 398 153 432 157
rect 862 289 896 323
rect 770 153 804 187
rect 954 249 988 255
rect 954 221 979 249
rect 979 221 988 249
rect 1142 221 1176 255
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
<< metal1 >>
rect 0 561 1656 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1656 561
rect 0 496 1656 527
rect 294 323 352 329
rect 294 289 306 323
rect 340 320 352 323
rect 850 323 908 329
rect 850 320 862 323
rect 340 292 862 320
rect 340 289 352 292
rect 294 283 352 289
rect 850 289 862 292
rect 896 289 908 323
rect 850 283 908 289
rect 942 255 1000 261
rect 942 221 954 255
rect 988 252 1000 255
rect 1130 255 1188 261
rect 1130 252 1142 255
rect 988 224 1142 252
rect 988 221 1000 224
rect 942 215 1000 221
rect 1130 221 1142 224
rect 1176 221 1188 255
rect 1130 215 1188 221
rect 386 187 444 193
rect 386 153 398 187
rect 432 184 444 187
rect 758 187 816 193
rect 758 184 770 187
rect 432 156 770 184
rect 432 153 444 156
rect 386 147 444 153
rect 758 153 770 156
rect 804 153 816 187
rect 758 147 816 153
rect 0 17 1656 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1656 17
rect 0 -48 1656 -17
<< labels >>
flabel locali s 30 289 64 323 0 FreeSans 200 0 0 0 SCE
port 3 nsew signal input
flabel locali s 954 221 988 255 0 FreeSans 200 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1326 425 1360 459 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1326 357 1360 391 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 214 357 248 391 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 1326 85 1360 119 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 214 289 248 323 0 FreeSans 200 0 0 0 GATE
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 SCE
port 3 nsew signal input
flabel locali s 1418 221 1452 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1510 425 1544 459 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1510 357 1544 391 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1510 289 1544 323 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1510 221 1544 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1602 221 1636 255 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel locali s 1510 153 1544 187 0 FreeSans 200 0 0 0 GCLK
port 8 nsew signal output
flabel metal1 s 30 -17 64 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 30 527 64 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
flabel nwell s 30 527 64 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel pwell s 30 -17 64 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 sdlclkp_4
rlabel locali s 1137 199 1213 265 1 CLK
port 1 nsew clock input
rlabel metal1 s 1130 252 1188 261 1 CLK
port 1 nsew clock input
rlabel metal1 s 1130 215 1188 224 1 CLK
port 1 nsew clock input
rlabel metal1 s 942 252 1000 261 1 CLK
port 1 nsew clock input
rlabel metal1 s 942 224 1188 252 1 CLK
port 1 nsew clock input
rlabel metal1 s 942 215 1000 224 1 CLK
port 1 nsew clock input
rlabel metal1 s 0 -48 1656 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1656 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1656 544
string GDS_END 444834
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 431426
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 8.280 0.000 
<< end >>
