magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 682 582
<< pwell >>
rect 1 21 643 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 174 47 204 177
rect 247 47 277 177
rect 435 47 465 177
rect 526 47 556 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 247 297 277 497
rect 435 297 465 497
rect 526 297 556 497
<< ndiff >>
rect 27 129 79 177
rect 27 95 35 129
rect 69 95 79 129
rect 27 47 79 95
rect 109 105 174 177
rect 109 71 119 105
rect 153 71 174 105
rect 109 47 174 71
rect 204 47 247 177
rect 277 101 329 177
rect 277 67 287 101
rect 321 67 329 101
rect 277 47 329 67
rect 383 101 435 177
rect 383 67 391 101
rect 425 67 435 101
rect 383 47 435 67
rect 465 47 526 177
rect 556 97 617 177
rect 556 63 566 97
rect 600 63 617 97
rect 556 47 617 63
<< pdiff >>
rect 27 477 79 497
rect 27 443 35 477
rect 69 443 79 477
rect 27 347 79 443
rect 27 313 35 347
rect 69 313 79 347
rect 27 297 79 313
rect 109 477 163 497
rect 109 443 119 477
rect 153 443 163 477
rect 109 409 163 443
rect 109 375 119 409
rect 153 375 163 409
rect 109 297 163 375
rect 193 409 247 497
rect 193 375 203 409
rect 237 375 247 409
rect 193 297 247 375
rect 277 485 329 497
rect 277 451 287 485
rect 321 451 329 485
rect 277 297 329 451
rect 383 477 435 497
rect 383 443 391 477
rect 425 443 435 477
rect 383 297 435 443
rect 465 477 526 497
rect 465 443 475 477
rect 509 443 526 477
rect 465 407 526 443
rect 465 373 475 407
rect 509 373 526 407
rect 465 297 526 373
rect 556 477 617 497
rect 556 443 575 477
rect 609 443 617 477
rect 556 409 617 443
rect 556 375 575 409
rect 609 375 617 409
rect 556 297 617 375
<< ndiffc >>
rect 35 95 69 129
rect 119 71 153 105
rect 287 67 321 101
rect 391 67 425 101
rect 566 63 600 97
<< pdiffc >>
rect 35 443 69 477
rect 35 313 69 347
rect 119 443 153 477
rect 119 375 153 409
rect 203 375 237 409
rect 287 451 321 485
rect 391 443 425 477
rect 475 443 509 477
rect 475 373 509 407
rect 575 443 609 477
rect 575 375 609 409
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 247 497 277 523
rect 435 497 465 523
rect 526 497 556 523
rect 79 265 109 297
rect 163 265 193 297
rect 247 265 277 297
rect 435 265 465 297
rect 526 265 556 297
rect 21 249 109 265
rect 21 215 33 249
rect 67 215 109 249
rect 21 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 249 306 265
rect 247 215 261 249
rect 295 215 306 249
rect 247 199 306 215
rect 395 249 465 265
rect 395 215 405 249
rect 439 215 465 249
rect 395 199 465 215
rect 507 249 561 265
rect 507 215 517 249
rect 551 215 561 249
rect 507 199 561 215
rect 79 177 109 199
rect 174 177 204 199
rect 247 177 277 199
rect 435 177 465 199
rect 526 177 556 199
rect 79 21 109 47
rect 174 21 204 47
rect 247 21 277 47
rect 435 21 465 47
rect 526 21 556 47
<< polycont >>
rect 33 215 67 249
rect 161 215 195 249
rect 261 215 295 249
rect 405 215 439 249
rect 517 215 551 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 35 477 69 493
rect 35 347 69 443
rect 103 485 337 493
rect 103 477 287 485
rect 103 443 119 477
rect 153 459 287 477
rect 271 451 287 459
rect 321 451 337 485
rect 375 477 441 527
rect 375 443 391 477
rect 425 443 441 477
rect 475 477 525 493
rect 509 443 525 477
rect 103 409 153 443
rect 103 375 119 409
rect 103 359 153 375
rect 203 409 248 425
rect 475 409 525 443
rect 237 407 525 409
rect 237 375 475 407
rect 203 373 475 375
rect 509 373 525 407
rect 559 477 625 527
rect 559 443 575 477
rect 609 443 625 477
rect 559 409 625 443
rect 559 375 575 409
rect 609 375 625 409
rect 203 367 525 373
rect 203 359 405 367
rect 430 325 627 333
rect 69 313 627 325
rect 35 299 627 313
rect 35 291 460 299
rect 17 249 87 257
rect 17 215 33 249
rect 67 215 87 249
rect 123 249 211 257
rect 123 215 161 249
rect 195 215 211 249
rect 245 249 339 257
rect 245 215 261 249
rect 295 215 339 249
rect 34 147 247 181
rect 34 129 69 147
rect 34 95 35 129
rect 34 51 69 95
rect 103 105 169 113
rect 103 71 119 105
rect 153 71 169 105
rect 103 17 169 71
rect 213 101 247 147
rect 283 135 339 215
rect 389 249 455 257
rect 389 215 405 249
rect 439 215 455 249
rect 494 249 551 265
rect 494 215 517 249
rect 389 135 440 215
rect 494 199 551 215
rect 585 165 627 299
rect 476 131 627 165
rect 476 101 516 131
rect 213 67 287 101
rect 321 67 391 101
rect 425 67 516 101
rect 213 51 516 67
rect 550 63 566 97
rect 600 63 616 97
rect 550 17 616 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
<< metal1 >>
rect 0 561 644 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 644 561
rect 0 496 644 527
rect 0 17 644 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 644 17
rect 0 -48 644 -17
<< labels >>
flabel locali s 586 153 620 187 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 586 289 620 323 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 586 221 620 255 0 FreeSans 200 0 0 0 Y
port 10 nsew signal output
flabel locali s 29 221 63 255 0 FreeSans 200 0 0 0 C1
port 5 nsew signal input
flabel locali s 397 221 431 255 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 494 221 528 255 0 FreeSans 200 0 0 0 A2
port 2 nsew signal input
flabel locali s 123 221 157 255 0 FreeSans 200 0 0 0 B2
port 4 nsew signal input
flabel locali s 305 221 339 255 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel locali s 397 153 431 187 0 FreeSans 200 0 0 0 A1
port 1 nsew signal input
flabel locali s 305 153 339 187 0 FreeSans 200 0 0 0 B1
port 3 nsew signal input
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 6 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 9 nsew power bidirectional abutment
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 8 nsew power bidirectional
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 7 nsew ground bidirectional
rlabel comment s 0 0 0 0 4 a221oi_1
rlabel metal1 s 0 -48 644 48 1 VGND
port 6 nsew ground bidirectional abutment
rlabel metal1 s 0 496 644 592 1 VPWR
port 9 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 644 544
string GDS_END 3590080
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3583510
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 16.100 0.000 
<< end >>
