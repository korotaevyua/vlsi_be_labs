magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 866 582
<< pwell >>
rect 1 21 808 203
rect 30 -17 64 21
<< locali >>
rect 119 265 166 410
rect 17 215 85 265
rect 119 215 211 265
rect 245 215 340 265
rect 469 325 519 493
rect 637 325 687 493
rect 469 291 811 325
rect 753 181 811 291
rect 461 147 811 181
rect 461 53 527 147
rect 629 53 695 147
<< obsli1 >>
rect 0 527 828 561
rect 17 459 253 493
rect 17 299 85 459
rect 200 333 253 459
rect 287 367 427 527
rect 200 299 418 333
rect 374 249 418 299
rect 553 359 603 527
rect 721 359 771 527
rect 374 215 719 249
rect 374 181 418 215
rect 17 145 418 181
rect 17 51 85 145
rect 119 17 153 111
rect 187 51 253 145
rect 287 17 427 111
rect 561 17 595 111
rect 729 17 763 111
rect 0 -17 828 17
<< metal1 >>
rect 0 496 828 592
rect 0 -48 828 48
<< labels >>
rlabel locali s 245 215 340 265 6 A
port 1 nsew signal input
rlabel locali s 119 215 211 265 6 B
port 2 nsew signal input
rlabel locali s 119 265 166 410 6 B
port 2 nsew signal input
rlabel locali s 17 215 85 265 6 C
port 3 nsew signal input
rlabel metal1 s 0 -48 828 48 8 VGND
port 4 nsew ground bidirectional abutment
rlabel pwell s 30 -17 64 21 6 VNB
port 5 nsew ground bidirectional
rlabel pwell s 1 21 808 203 6 VNB
port 5 nsew ground bidirectional
rlabel nwell s -38 261 866 582 6 VPB
port 6 nsew power bidirectional
rlabel metal1 s 0 496 828 592 6 VPWR
port 7 nsew power bidirectional abutment
rlabel locali s 629 53 695 147 6 X
port 8 nsew signal output
rlabel locali s 461 53 527 147 6 X
port 8 nsew signal output
rlabel locali s 461 147 811 181 6 X
port 8 nsew signal output
rlabel locali s 753 181 811 291 6 X
port 8 nsew signal output
rlabel locali s 469 291 811 325 6 X
port 8 nsew signal output
rlabel locali s 637 325 687 493 6 X
port 8 nsew signal output
rlabel locali s 469 325 519 493 6 X
port 8 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 828 544
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1029624
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1022566
<< end >>
