magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 130 827
rect 384 261 596 827
rect 850 261 1481 827
<< pwell >>
rect 3 893 89 1050
rect 511 885 1111 1067
rect 1383 893 1469 1050
rect 3 38 89 195
rect 601 192 1425 203
rect 398 56 1425 192
rect 601 21 1425 56
<< locali >>
rect 594 214 658 308
rect 1072 282 1127 474
rect 1256 282 1311 474
rect 1072 217 1311 282
rect 1072 196 1127 217
rect 1067 51 1127 196
rect 1267 51 1311 217
<< obsli1 >>
rect 0 1071 1472 1105
rect 17 926 75 1071
rect 529 903 581 1071
rect 615 865 681 1037
rect 715 903 753 1071
rect 787 865 853 1037
rect 889 903 991 1071
rect 1027 964 1097 1032
rect 1027 892 1139 964
rect 1397 926 1455 1071
rect 1027 881 1153 892
rect 615 853 853 865
rect 1072 871 1153 881
rect 629 831 839 853
rect 17 597 75 794
rect 0 527 378 561
rect 412 532 562 750
rect 412 467 478 532
rect 612 474 678 793
rect 804 762 838 831
rect 1072 825 1217 871
rect 882 728 944 748
rect 736 694 944 728
rect 736 515 770 694
rect 804 583 838 660
rect 878 617 944 694
rect 804 549 928 583
rect 736 481 838 515
rect 276 413 478 467
rect 412 327 478 413
rect 512 426 678 474
rect 17 17 75 162
rect 404 17 470 179
rect 512 75 560 426
rect 804 196 838 481
rect 894 325 928 549
rect 978 561 1024 748
rect 1072 614 1110 825
rect 1397 597 1455 791
rect 978 527 1472 561
rect 978 325 1024 527
rect 1181 322 1215 527
rect 1351 322 1387 527
rect 623 17 689 180
rect 723 146 933 196
rect 723 51 761 146
rect 795 17 861 112
rect 895 51 933 146
rect 967 17 1033 180
rect 1165 17 1231 169
rect 1351 17 1401 185
rect 0 -17 1472 17
<< metal1 >>
rect 0 1040 1472 1136
rect 16 728 74 737
rect 1386 728 1444 737
rect 14 700 1458 728
rect 16 691 74 700
rect 1386 691 1444 700
rect 0 496 1472 592
rect 272 456 474 463
rect 14 428 1458 456
rect 272 417 474 428
rect 0 -48 1472 48
<< labels >>
rlabel locali s 594 214 658 308 6 A
port 1 nsew signal input
rlabel metal1 s 0 1040 1472 1136 6 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 1383 893 1469 1050 6 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 3 893 89 1050 6 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 0 -48 1472 48 8 VGND
port 2 nsew ground bidirectional abutment
rlabel pwell s 3 38 89 195 6 VGND
port 2 nsew ground bidirectional abutment
rlabel metal1 s 1386 691 1444 700 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 16 691 74 700 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 14 700 1458 728 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 1386 728 1444 737 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 16 728 74 737 6 VPB
port 3 nsew power bidirectional
rlabel nwell s 850 261 1481 827 6 VPB
port 3 nsew power bidirectional
rlabel nwell s -38 261 130 827 6 VPB
port 3 nsew power bidirectional
rlabel metal1 s 272 417 474 428 6 VPWRIN
port 4 nsew power bidirectional abutment
rlabel metal1 s 14 428 1458 456 6 VPWRIN
port 4 nsew power bidirectional abutment
rlabel metal1 s 272 456 474 463 6 VPWRIN
port 4 nsew power bidirectional abutment
rlabel nwell s 384 261 596 827 6 VPWRIN
port 4 nsew power bidirectional abutment
rlabel metal1 s 0 496 1472 592 6 VPWR
port 5 nsew power bidirectional abutment
rlabel locali s 1267 51 1311 217 6 X
port 6 nsew signal output
rlabel locali s 1067 51 1127 196 6 X
port 6 nsew signal output
rlabel locali s 1072 196 1127 217 6 X
port 6 nsew signal output
rlabel locali s 1072 217 1311 282 6 X
port 6 nsew signal output
rlabel locali s 1256 282 1311 474 6 X
port 6 nsew signal output
rlabel locali s 1072 282 1127 474 6 X
port 6 nsew signal output
<< properties >>
string FIXED_BBOX 0 0 1472 1088
string LEFclass CORE WELLTAP
string LEFsite unithd
string LEFsymmetry X Y R90
string LEFview TRUE
string GDS_END 1567436
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1552930
<< end >>
