magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 1234 582
<< pwell >>
rect 16 21 1183 203
rect 29 -17 63 21
<< scnmos >>
rect 119 47 149 177
rect 205 47 235 177
rect 291 47 321 177
rect 377 47 407 177
rect 463 47 493 177
rect 655 47 685 177
rect 739 47 769 177
rect 831 47 861 177
rect 907 47 937 177
rect 991 47 1021 177
rect 1075 47 1105 177
<< scpmoshvt >>
rect 119 297 149 497
rect 205 297 235 497
rect 291 297 321 497
rect 377 297 407 497
rect 463 297 493 497
rect 655 297 685 497
rect 739 297 769 497
rect 823 297 853 497
rect 907 297 937 497
rect 991 297 1021 497
rect 1075 297 1105 497
<< ndiff >>
rect 42 157 119 177
rect 42 123 58 157
rect 92 123 119 157
rect 42 89 119 123
rect 42 55 58 89
rect 92 55 119 89
rect 42 47 119 55
rect 149 89 205 177
rect 149 55 160 89
rect 194 55 205 89
rect 149 47 205 55
rect 235 157 291 177
rect 235 123 246 157
rect 280 123 291 157
rect 235 47 291 123
rect 321 89 377 177
rect 321 55 332 89
rect 366 55 377 89
rect 321 47 377 55
rect 407 157 463 177
rect 407 123 418 157
rect 452 123 463 157
rect 407 47 463 123
rect 493 89 655 177
rect 493 55 526 89
rect 560 55 607 89
rect 641 55 655 89
rect 493 47 655 55
rect 685 169 739 177
rect 685 135 695 169
rect 729 135 739 169
rect 685 101 739 135
rect 685 67 695 101
rect 729 67 739 101
rect 685 47 739 67
rect 769 89 831 177
rect 769 55 787 89
rect 821 55 831 89
rect 769 47 831 55
rect 861 47 907 177
rect 937 131 991 177
rect 937 97 947 131
rect 981 97 991 131
rect 937 47 991 97
rect 1021 47 1075 177
rect 1105 161 1157 177
rect 1105 127 1115 161
rect 1149 127 1157 161
rect 1105 93 1157 127
rect 1105 59 1115 93
rect 1149 59 1157 93
rect 1105 47 1157 59
<< pdiff >>
rect 66 477 119 497
rect 66 443 74 477
rect 108 443 119 477
rect 66 409 119 443
rect 66 375 74 409
rect 108 375 119 409
rect 66 297 119 375
rect 149 489 205 497
rect 149 455 160 489
rect 194 455 205 489
rect 149 297 205 455
rect 235 353 291 497
rect 235 319 246 353
rect 280 319 291 353
rect 235 297 291 319
rect 321 489 377 497
rect 321 455 332 489
rect 366 455 377 489
rect 321 297 377 455
rect 407 353 463 497
rect 407 319 418 353
rect 452 319 463 353
rect 407 297 463 319
rect 493 489 549 497
rect 493 455 503 489
rect 537 455 549 489
rect 493 297 549 455
rect 603 459 655 497
rect 603 425 611 459
rect 645 425 655 459
rect 603 389 655 425
rect 603 355 611 389
rect 645 355 655 389
rect 603 297 655 355
rect 685 341 739 497
rect 685 307 695 341
rect 729 307 739 341
rect 685 297 739 307
rect 769 428 823 497
rect 769 394 779 428
rect 813 394 823 428
rect 769 339 823 394
rect 769 305 779 339
rect 813 305 823 339
rect 769 297 823 305
rect 853 489 907 497
rect 853 455 863 489
rect 897 455 907 489
rect 853 297 907 455
rect 937 421 991 497
rect 937 387 947 421
rect 981 387 991 421
rect 937 297 991 387
rect 1021 489 1075 497
rect 1021 455 1031 489
rect 1065 455 1075 489
rect 1021 297 1075 455
rect 1105 419 1157 497
rect 1105 385 1115 419
rect 1149 385 1157 419
rect 1105 343 1157 385
rect 1105 309 1115 343
rect 1149 309 1157 343
rect 1105 297 1157 309
<< ndiffc >>
rect 58 123 92 157
rect 58 55 92 89
rect 160 55 194 89
rect 246 123 280 157
rect 332 55 366 89
rect 418 123 452 157
rect 526 55 560 89
rect 607 55 641 89
rect 695 135 729 169
rect 695 67 729 101
rect 787 55 821 89
rect 947 97 981 131
rect 1115 127 1149 161
rect 1115 59 1149 93
<< pdiffc >>
rect 74 443 108 477
rect 74 375 108 409
rect 160 455 194 489
rect 246 319 280 353
rect 332 455 366 489
rect 418 319 452 353
rect 503 455 537 489
rect 611 425 645 459
rect 611 355 645 389
rect 695 307 729 341
rect 779 394 813 428
rect 779 305 813 339
rect 863 455 897 489
rect 947 387 981 421
rect 1031 455 1065 489
rect 1115 385 1149 419
rect 1115 309 1149 343
<< poly >>
rect 119 497 149 523
rect 205 497 235 523
rect 291 497 321 523
rect 377 497 407 523
rect 463 497 493 523
rect 655 497 685 523
rect 739 497 769 523
rect 823 497 853 523
rect 907 497 937 523
rect 991 497 1021 523
rect 1075 497 1105 523
rect 119 265 149 297
rect 205 265 235 297
rect 291 265 321 297
rect 377 265 407 297
rect 463 265 493 297
rect 655 265 685 297
rect 739 265 769 297
rect 823 265 853 297
rect 907 265 937 297
rect 991 265 1021 297
rect 106 249 160 265
rect 106 215 116 249
rect 150 215 160 249
rect 106 199 160 215
rect 205 249 516 265
rect 205 215 336 249
rect 370 215 404 249
rect 438 215 472 249
rect 506 215 516 249
rect 205 199 516 215
rect 617 249 769 265
rect 617 215 627 249
rect 661 215 769 249
rect 617 199 769 215
rect 811 249 865 265
rect 811 215 821 249
rect 855 215 865 249
rect 811 199 865 215
rect 907 249 1021 265
rect 907 215 941 249
rect 975 215 1021 249
rect 907 199 1021 215
rect 119 177 149 199
rect 205 177 235 199
rect 291 177 321 199
rect 377 177 407 199
rect 463 177 493 199
rect 655 177 685 199
rect 739 177 769 199
rect 831 177 861 199
rect 907 177 937 199
rect 991 177 1021 199
rect 1075 265 1105 297
rect 1075 249 1129 265
rect 1075 215 1085 249
rect 1119 215 1129 249
rect 1075 199 1129 215
rect 1075 177 1105 199
rect 119 21 149 47
rect 205 21 235 47
rect 291 21 321 47
rect 377 21 407 47
rect 463 21 493 47
rect 655 21 685 47
rect 739 21 769 47
rect 831 21 861 47
rect 907 21 937 47
rect 991 21 1021 47
rect 1075 21 1105 47
<< polycont >>
rect 116 215 150 249
rect 336 215 370 249
rect 404 215 438 249
rect 472 215 506 249
rect 627 215 661 249
rect 821 215 855 249
rect 941 215 975 249
rect 1085 215 1119 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 21 477 110 493
rect 21 443 74 477
rect 108 443 110 477
rect 144 489 210 527
rect 144 455 160 489
rect 194 455 210 489
rect 316 489 382 527
rect 316 455 332 489
rect 366 455 382 489
rect 487 489 554 527
rect 487 455 503 489
rect 537 455 554 489
rect 847 489 913 527
rect 611 459 813 476
rect 21 421 110 443
rect 645 442 813 459
rect 847 455 863 489
rect 897 455 913 489
rect 1015 489 1081 527
rect 1015 455 1031 489
rect 1065 455 1081 489
rect 21 409 574 421
rect 21 375 74 409
rect 108 387 574 409
rect 108 375 113 387
rect 21 359 113 375
rect 21 168 66 359
rect 100 249 166 325
rect 100 215 116 249
rect 150 215 166 249
rect 100 202 166 215
rect 200 319 246 353
rect 280 319 418 353
rect 452 319 482 353
rect 21 157 108 168
rect 21 123 58 157
rect 92 123 108 157
rect 200 157 247 319
rect 540 305 574 387
rect 611 389 645 425
rect 777 428 813 442
rect 777 394 779 428
rect 813 394 947 421
rect 777 387 947 394
rect 981 419 1165 421
rect 981 387 1115 419
rect 611 339 645 355
rect 695 341 729 361
rect 540 271 661 305
rect 281 249 506 265
rect 281 215 336 249
rect 370 215 404 249
rect 438 215 472 249
rect 599 249 661 271
rect 506 215 562 237
rect 281 199 562 215
rect 599 215 627 249
rect 599 199 661 215
rect 528 160 562 199
rect 695 169 729 307
rect 777 339 813 387
rect 1114 385 1115 387
rect 1149 385 1165 419
rect 777 305 779 339
rect 777 289 813 305
rect 849 319 1078 353
rect 849 255 884 319
rect 805 249 884 255
rect 805 215 821 249
rect 855 215 884 249
rect 805 202 884 215
rect 918 249 991 272
rect 918 215 941 249
rect 975 215 991 249
rect 918 202 991 215
rect 1044 258 1078 319
rect 1114 343 1165 385
rect 1114 309 1115 343
rect 1149 309 1165 343
rect 1114 292 1165 309
rect 1044 249 1140 258
rect 1044 215 1085 249
rect 1119 215 1140 249
rect 1044 211 1140 215
rect 528 157 602 160
rect 200 123 246 157
rect 280 123 418 157
rect 452 123 468 157
rect 528 135 695 157
rect 729 135 993 168
rect 528 134 993 135
rect 528 123 729 134
rect 21 89 108 123
rect 695 101 729 123
rect 21 55 58 89
rect 92 55 108 89
rect 21 51 108 55
rect 142 55 160 89
rect 194 55 210 89
rect 142 17 210 55
rect 316 55 332 89
rect 366 55 382 89
rect 316 17 382 55
rect 503 55 526 89
rect 560 55 607 89
rect 641 55 657 89
rect 503 17 657 55
rect 937 131 993 134
rect 937 97 947 131
rect 981 97 993 131
rect 695 51 729 67
rect 771 55 787 89
rect 821 55 837 89
rect 937 81 993 97
rect 1109 161 1165 177
rect 1109 127 1115 161
rect 1149 127 1165 161
rect 1109 93 1165 127
rect 771 17 837 55
rect 1109 59 1115 93
rect 1149 59 1165 93
rect 1109 17 1165 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
<< metal1 >>
rect 0 561 1196 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1196 561
rect 0 496 1196 527
rect 0 17 1196 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1196 17
rect 0 -48 1196 -17
<< labels >>
flabel locali s 121 221 155 255 0 FreeSans 340 0 0 0 B1_N
port 3 nsew signal input
flabel locali s 1044 289 1078 323 0 FreeSans 340 0 0 0 A2
port 2 nsew signal input
flabel locali s 952 221 986 255 0 FreeSans 340 0 0 0 A1
port 1 nsew signal input
flabel locali s 213 289 247 323 0 FreeSans 340 0 0 0 X
port 8 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 5 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 6 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 4 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 7 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 a21bo_4
rlabel metal1 s 0 -48 1196 48 1 VGND
port 4 nsew ground bidirectional abutment
rlabel metal1 s 0 496 1196 592 1 VPWR
port 7 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 1196 544
string GDS_END 3982802
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 3974554
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 29.900 0.000 
<< end >>
