magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 2430 582
<< pwell >>
rect 1173 157 1355 201
rect 1661 157 2390 203
rect 1 145 825 157
rect 1027 145 2390 157
rect 1 21 2390 145
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 131
rect 163 47 193 131
rect 355 47 385 131
rect 457 47 487 131
rect 535 47 565 131
rect 631 47 661 131
rect 707 47 737 131
rect 909 47 939 119
rect 1005 47 1035 119
rect 1103 47 1133 131
rect 1249 47 1279 175
rect 1350 47 1380 119
rect 1453 47 1483 119
rect 1548 47 1578 131
rect 1739 47 1769 177
rect 1827 47 1857 177
rect 1911 47 1941 177
rect 2101 47 2131 131
rect 2198 47 2228 177
rect 2282 47 2312 177
<< scpmoshvt >>
rect 80 363 110 491
rect 164 363 194 491
rect 352 369 382 497
rect 436 369 466 497
rect 530 369 560 497
rect 614 369 644 497
rect 707 369 737 497
rect 908 413 938 497
rect 1001 413 1031 497
rect 1097 413 1127 497
rect 1229 347 1259 497
rect 1324 413 1354 497
rect 1408 413 1438 497
rect 1525 413 1555 497
rect 1739 297 1769 497
rect 1827 297 1857 497
rect 1911 297 1941 497
rect 2101 369 2131 497
rect 2198 297 2228 497
rect 2282 297 2312 497
<< ndiff >>
rect 27 119 79 131
rect 27 85 35 119
rect 69 85 79 119
rect 27 47 79 85
rect 109 93 163 131
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 119 245 131
rect 193 85 203 119
rect 237 85 245 119
rect 193 47 245 85
rect 299 89 355 131
rect 299 55 311 89
rect 345 55 355 89
rect 299 47 355 55
rect 385 89 457 131
rect 385 55 411 89
rect 445 55 457 89
rect 385 47 457 55
rect 487 47 535 131
rect 565 89 631 131
rect 565 55 586 89
rect 620 55 631 89
rect 565 47 631 55
rect 661 47 707 131
rect 737 89 799 131
rect 1199 131 1249 175
rect 1053 119 1103 131
rect 737 55 753 89
rect 787 55 799 89
rect 737 47 799 55
rect 853 107 909 119
rect 853 73 861 107
rect 895 73 909 107
rect 853 47 909 73
rect 939 107 1005 119
rect 939 73 961 107
rect 995 73 1005 107
rect 939 47 1005 73
rect 1035 47 1103 119
rect 1133 101 1249 131
rect 1133 67 1177 101
rect 1211 67 1249 101
rect 1133 47 1249 67
rect 1279 119 1329 175
rect 1687 162 1739 177
rect 1498 119 1548 131
rect 1279 107 1350 119
rect 1279 73 1295 107
rect 1329 73 1350 107
rect 1279 47 1350 73
rect 1380 107 1453 119
rect 1380 73 1407 107
rect 1441 73 1453 107
rect 1380 47 1453 73
rect 1483 47 1548 119
rect 1578 107 1630 131
rect 1578 73 1588 107
rect 1622 73 1630 107
rect 1578 47 1630 73
rect 1687 128 1695 162
rect 1729 128 1739 162
rect 1687 94 1739 128
rect 1687 60 1695 94
rect 1729 60 1739 94
rect 1687 47 1739 60
rect 1769 123 1827 177
rect 1769 89 1781 123
rect 1815 89 1827 123
rect 1769 47 1827 89
rect 1857 157 1911 177
rect 1857 123 1867 157
rect 1901 123 1911 157
rect 1857 89 1911 123
rect 1857 55 1867 89
rect 1901 55 1911 89
rect 1857 47 1911 55
rect 1941 122 1995 177
rect 2146 161 2198 177
rect 2146 131 2154 161
rect 1941 88 1953 122
rect 1987 88 1995 122
rect 1941 47 1995 88
rect 2049 119 2101 131
rect 2049 85 2057 119
rect 2091 85 2101 119
rect 2049 47 2101 85
rect 2131 127 2154 131
rect 2188 127 2198 161
rect 2131 93 2198 127
rect 2131 59 2154 93
rect 2188 59 2198 93
rect 2131 47 2198 59
rect 2228 143 2282 177
rect 2228 109 2238 143
rect 2272 109 2282 143
rect 2228 47 2282 109
rect 2312 161 2364 177
rect 2312 127 2322 161
rect 2356 127 2364 161
rect 2312 93 2364 127
rect 2312 59 2322 93
rect 2356 59 2364 93
rect 2312 47 2364 59
<< pdiff >>
rect 28 477 80 491
rect 28 443 36 477
rect 70 443 80 477
rect 28 409 80 443
rect 28 375 36 409
rect 70 375 80 409
rect 28 363 80 375
rect 110 461 164 491
rect 110 427 120 461
rect 154 427 164 461
rect 110 363 164 427
rect 194 477 246 491
rect 194 443 204 477
rect 238 443 246 477
rect 194 409 246 443
rect 194 375 204 409
rect 238 375 246 409
rect 194 363 246 375
rect 300 452 352 497
rect 300 418 308 452
rect 342 418 352 452
rect 300 369 352 418
rect 382 483 436 497
rect 382 449 392 483
rect 426 449 436 483
rect 382 369 436 449
rect 466 369 530 497
rect 560 483 614 497
rect 560 449 570 483
rect 604 449 614 483
rect 560 369 614 449
rect 644 369 707 497
rect 737 483 794 497
rect 737 449 752 483
rect 786 449 794 483
rect 737 369 794 449
rect 855 472 908 497
rect 855 438 863 472
rect 897 438 908 472
rect 855 413 908 438
rect 938 472 1001 497
rect 938 438 953 472
rect 987 438 1001 472
rect 938 413 1001 438
rect 1031 413 1097 497
rect 1127 485 1229 497
rect 1127 451 1185 485
rect 1219 451 1229 485
rect 1127 417 1229 451
rect 1127 413 1185 417
rect 1142 383 1185 413
rect 1219 383 1229 417
rect 1142 347 1229 383
rect 1259 477 1324 497
rect 1259 443 1269 477
rect 1303 443 1324 477
rect 1259 413 1324 443
rect 1354 467 1408 497
rect 1354 433 1364 467
rect 1398 433 1408 467
rect 1354 413 1408 433
rect 1438 413 1525 497
rect 1555 477 1630 497
rect 1555 443 1587 477
rect 1621 443 1630 477
rect 1555 413 1630 443
rect 1687 485 1739 497
rect 1687 451 1695 485
rect 1729 451 1739 485
rect 1687 417 1739 451
rect 1259 347 1309 413
rect 1687 383 1695 417
rect 1729 383 1739 417
rect 1687 349 1739 383
rect 1687 315 1695 349
rect 1729 315 1739 349
rect 1687 297 1739 315
rect 1769 455 1827 497
rect 1769 421 1781 455
rect 1815 421 1827 455
rect 1769 375 1827 421
rect 1769 341 1781 375
rect 1815 341 1827 375
rect 1769 297 1827 341
rect 1857 479 1911 497
rect 1857 445 1867 479
rect 1901 445 1911 479
rect 1857 411 1911 445
rect 1857 377 1867 411
rect 1901 377 1911 411
rect 1857 343 1911 377
rect 1857 309 1867 343
rect 1901 309 1911 343
rect 1857 297 1911 309
rect 1941 485 1995 497
rect 1941 451 1953 485
rect 1987 451 1995 485
rect 1941 373 1995 451
rect 1941 339 1953 373
rect 1987 339 1995 373
rect 2049 485 2101 497
rect 2049 451 2057 485
rect 2091 451 2101 485
rect 2049 417 2101 451
rect 2049 383 2057 417
rect 2091 383 2101 417
rect 2049 369 2101 383
rect 2131 485 2198 497
rect 2131 451 2154 485
rect 2188 451 2198 485
rect 2131 417 2198 451
rect 2131 383 2154 417
rect 2188 383 2198 417
rect 2131 369 2198 383
rect 1941 297 1995 339
rect 2146 349 2198 369
rect 2146 315 2154 349
rect 2188 315 2198 349
rect 2146 297 2198 315
rect 2228 449 2282 497
rect 2228 415 2238 449
rect 2272 415 2282 449
rect 2228 381 2282 415
rect 2228 347 2238 381
rect 2272 347 2282 381
rect 2228 297 2282 347
rect 2312 485 2364 497
rect 2312 451 2322 485
rect 2356 451 2364 485
rect 2312 417 2364 451
rect 2312 383 2322 417
rect 2356 383 2364 417
rect 2312 349 2364 383
rect 2312 315 2322 349
rect 2356 315 2364 349
rect 2312 297 2364 315
<< ndiffc >>
rect 35 85 69 119
rect 119 59 153 93
rect 203 85 237 119
rect 311 55 345 89
rect 411 55 445 89
rect 586 55 620 89
rect 753 55 787 89
rect 861 73 895 107
rect 961 73 995 107
rect 1177 67 1211 101
rect 1295 73 1329 107
rect 1407 73 1441 107
rect 1588 73 1622 107
rect 1695 128 1729 162
rect 1695 60 1729 94
rect 1781 89 1815 123
rect 1867 123 1901 157
rect 1867 55 1901 89
rect 1953 88 1987 122
rect 2057 85 2091 119
rect 2154 127 2188 161
rect 2154 59 2188 93
rect 2238 109 2272 143
rect 2322 127 2356 161
rect 2322 59 2356 93
<< pdiffc >>
rect 36 443 70 477
rect 36 375 70 409
rect 120 427 154 461
rect 204 443 238 477
rect 204 375 238 409
rect 308 418 342 452
rect 392 449 426 483
rect 570 449 604 483
rect 752 449 786 483
rect 863 438 897 472
rect 953 438 987 472
rect 1185 451 1219 485
rect 1185 383 1219 417
rect 1269 443 1303 477
rect 1364 433 1398 467
rect 1587 443 1621 477
rect 1695 451 1729 485
rect 1695 383 1729 417
rect 1695 315 1729 349
rect 1781 421 1815 455
rect 1781 341 1815 375
rect 1867 445 1901 479
rect 1867 377 1901 411
rect 1867 309 1901 343
rect 1953 451 1987 485
rect 1953 339 1987 373
rect 2057 451 2091 485
rect 2057 383 2091 417
rect 2154 451 2188 485
rect 2154 383 2188 417
rect 2154 315 2188 349
rect 2238 415 2272 449
rect 2238 347 2272 381
rect 2322 451 2356 485
rect 2322 383 2356 417
rect 2322 315 2356 349
<< poly >>
rect 80 491 110 517
rect 164 491 194 517
rect 352 497 382 523
rect 436 497 466 523
rect 530 497 560 523
rect 614 497 644 523
rect 707 497 737 523
rect 908 497 938 523
rect 1001 497 1031 523
rect 1097 497 1127 523
rect 1229 497 1259 523
rect 1324 497 1354 523
rect 1408 497 1438 523
rect 1525 497 1555 523
rect 1739 497 1769 523
rect 1827 497 1857 523
rect 1911 497 1941 523
rect 2101 497 2131 523
rect 2198 497 2228 523
rect 2282 497 2312 523
rect 908 375 938 413
rect 1001 381 1031 413
rect 80 348 110 363
rect 47 318 110 348
rect 47 265 77 318
rect 164 274 194 363
rect 352 331 382 369
rect 436 331 466 369
rect 530 337 560 369
rect 614 337 644 369
rect 340 321 466 331
rect 340 287 356 321
rect 390 301 466 321
rect 515 321 569 337
rect 390 287 406 301
rect 340 277 406 287
rect 515 287 525 321
rect 559 287 569 321
rect 23 249 77 265
rect 23 215 33 249
rect 67 215 77 249
rect 119 264 194 274
rect 119 230 135 264
rect 169 230 194 264
rect 119 220 194 230
rect 23 199 77 215
rect 47 176 77 199
rect 47 146 109 176
rect 79 131 109 146
rect 163 131 193 220
rect 355 131 385 277
rect 515 271 569 287
rect 611 321 665 337
rect 611 287 621 321
rect 655 287 665 321
rect 611 271 665 287
rect 707 304 737 369
rect 893 365 959 375
rect 893 331 909 365
rect 943 331 959 365
rect 893 321 959 331
rect 1001 365 1055 381
rect 1001 331 1011 365
rect 1045 331 1055 365
rect 1001 315 1055 331
rect 707 288 761 304
rect 427 225 493 235
rect 427 191 443 225
rect 477 191 493 225
rect 427 181 493 191
rect 457 131 487 181
rect 535 131 565 271
rect 707 254 717 288
rect 751 254 761 288
rect 1001 279 1031 315
rect 707 238 761 254
rect 909 249 1031 279
rect 607 207 661 223
rect 607 173 617 207
rect 651 173 661 207
rect 607 157 661 173
rect 631 131 661 157
rect 707 131 737 238
rect 909 119 939 249
rect 1097 213 1127 413
rect 1229 309 1259 347
rect 1324 315 1354 413
rect 1408 375 1438 413
rect 1525 381 1555 413
rect 1407 365 1473 375
rect 1407 331 1423 365
rect 1457 331 1473 365
rect 1407 321 1473 331
rect 1525 365 1603 381
rect 1525 331 1559 365
rect 1593 331 1603 365
rect 1525 315 1603 331
rect 1169 299 1259 309
rect 1169 265 1185 299
rect 1219 265 1259 299
rect 1169 255 1259 265
rect 1229 220 1259 255
rect 1311 299 1365 315
rect 1311 265 1321 299
rect 1355 279 1365 299
rect 1355 265 1483 279
rect 1311 249 1483 265
rect 981 191 1035 207
rect 981 157 991 191
rect 1025 157 1035 191
rect 1097 203 1177 213
rect 1097 183 1127 203
rect 981 141 1035 157
rect 1005 119 1035 141
rect 1103 169 1127 183
rect 1161 169 1177 203
rect 1229 190 1279 220
rect 1249 175 1279 190
rect 1350 191 1411 207
rect 1103 159 1177 169
rect 1103 131 1133 159
rect 1350 157 1367 191
rect 1401 157 1411 191
rect 1350 141 1411 157
rect 1350 119 1380 141
rect 1453 119 1483 249
rect 1548 131 1578 315
rect 2101 333 2131 369
rect 2090 303 2131 333
rect 1739 265 1769 297
rect 1827 265 1857 297
rect 1911 265 1941 297
rect 2090 265 2120 303
rect 2198 265 2228 297
rect 2282 265 2312 297
rect 1630 249 1769 265
rect 1630 215 1640 249
rect 1674 215 1769 249
rect 1630 199 1769 215
rect 1811 249 2120 265
rect 1811 215 1821 249
rect 1855 215 2120 249
rect 1811 199 2120 215
rect 2169 249 2312 265
rect 2169 215 2179 249
rect 2213 215 2312 249
rect 2169 199 2312 215
rect 1739 177 1769 199
rect 1827 177 1857 199
rect 1911 177 1941 199
rect 2090 176 2120 199
rect 2198 177 2228 199
rect 2282 177 2312 199
rect 2090 146 2131 176
rect 2101 131 2131 146
rect 79 21 109 47
rect 163 21 193 47
rect 355 21 385 47
rect 457 21 487 47
rect 535 21 565 47
rect 631 21 661 47
rect 707 21 737 47
rect 909 21 939 47
rect 1005 21 1035 47
rect 1103 21 1133 47
rect 1249 21 1279 47
rect 1350 21 1380 47
rect 1453 21 1483 47
rect 1548 21 1578 47
rect 1739 21 1769 47
rect 1827 21 1857 47
rect 1911 21 1941 47
rect 2101 21 2131 47
rect 2198 21 2228 47
rect 2282 21 2312 47
<< polycont >>
rect 356 287 390 321
rect 525 287 559 321
rect 33 215 67 249
rect 135 230 169 264
rect 621 287 655 321
rect 909 331 943 365
rect 1011 331 1045 365
rect 443 191 477 225
rect 717 254 751 288
rect 617 173 651 207
rect 1423 331 1457 365
rect 1559 331 1593 365
rect 1185 265 1219 299
rect 1321 265 1355 299
rect 991 157 1025 191
rect 1127 169 1161 203
rect 1367 157 1401 191
rect 1640 215 1674 249
rect 1821 215 1855 249
rect 2179 215 2213 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 36 477 70 493
rect 36 409 70 443
rect 104 461 170 527
rect 104 427 120 461
rect 154 427 170 461
rect 204 477 249 493
rect 238 443 249 477
rect 204 409 249 443
rect 70 391 169 393
rect 70 375 129 391
rect 36 359 129 375
rect 123 357 129 359
rect 163 357 169 391
rect 19 249 89 325
rect 19 215 33 249
rect 67 215 89 249
rect 19 195 89 215
rect 123 264 169 357
rect 123 230 135 264
rect 123 194 169 230
rect 238 375 249 409
rect 123 161 162 194
rect 35 127 162 161
rect 204 187 249 375
rect 204 153 210 187
rect 244 153 249 187
rect 204 143 249 153
rect 35 119 69 127
rect 203 119 249 143
rect 35 69 69 85
rect 103 59 119 93
rect 153 59 169 93
rect 237 85 249 119
rect 203 69 249 85
rect 287 452 342 489
rect 287 418 308 452
rect 376 483 442 527
rect 752 483 786 527
rect 376 449 392 483
rect 426 449 442 483
rect 539 449 570 483
rect 604 449 718 483
rect 287 415 342 418
rect 287 372 650 415
rect 287 89 321 372
rect 356 321 390 337
rect 356 157 390 287
rect 424 225 458 372
rect 616 337 650 372
rect 684 399 718 449
rect 752 433 786 449
rect 841 472 897 488
rect 1185 485 1219 527
rect 841 438 863 472
rect 937 438 953 472
rect 987 438 1151 472
rect 841 413 897 438
rect 841 399 875 413
rect 684 365 875 399
rect 995 391 1083 402
rect 492 321 559 337
rect 492 287 525 321
rect 492 271 559 287
rect 616 321 655 337
rect 616 287 621 321
rect 616 271 655 287
rect 707 288 807 331
rect 707 254 717 288
rect 751 254 807 288
rect 424 191 443 225
rect 477 191 493 225
rect 617 207 651 223
rect 707 207 807 254
rect 841 173 875 365
rect 617 157 651 173
rect 356 123 651 157
rect 685 139 875 173
rect 909 365 957 381
rect 943 331 957 365
rect 995 365 1041 391
rect 995 331 1011 365
rect 1075 357 1083 391
rect 1045 331 1083 357
rect 909 207 957 331
rect 1117 315 1151 438
rect 1185 417 1219 451
rect 1185 367 1219 383
rect 1253 477 1303 493
rect 1253 443 1269 477
rect 1561 477 1622 527
rect 1253 427 1303 443
rect 1348 433 1364 467
rect 1398 433 1525 467
rect 1117 299 1219 315
rect 1117 297 1185 299
rect 1059 265 1185 297
rect 1059 263 1219 265
rect 909 191 1025 207
rect 909 187 991 191
rect 909 153 949 187
rect 983 157 991 187
rect 983 153 1025 157
rect 909 141 1025 153
rect 103 17 169 59
rect 287 55 311 89
rect 345 55 361 89
rect 395 55 411 89
rect 445 55 461 89
rect 495 61 530 123
rect 685 89 719 139
rect 841 107 875 139
rect 1059 107 1093 263
rect 1185 249 1219 263
rect 1127 213 1161 219
rect 1253 213 1287 427
rect 1321 391 1359 393
rect 1321 357 1325 391
rect 1321 299 1359 357
rect 1355 265 1359 299
rect 1321 249 1359 265
rect 1393 365 1457 381
rect 1393 331 1423 365
rect 1393 315 1457 331
rect 1127 203 1287 213
rect 1393 207 1431 315
rect 1491 281 1525 433
rect 1561 443 1587 477
rect 1621 443 1622 477
rect 1561 427 1622 443
rect 1679 485 1745 491
rect 1679 451 1695 485
rect 1729 451 1745 485
rect 1679 417 1745 451
rect 1679 383 1695 417
rect 1729 383 1745 417
rect 1679 381 1745 383
rect 1559 365 1745 381
rect 1593 349 1745 365
rect 1593 331 1695 349
rect 1559 315 1695 331
rect 1729 315 1745 349
rect 1779 455 1815 527
rect 1779 421 1781 455
rect 1779 375 1815 421
rect 1779 341 1781 375
rect 1779 325 1815 341
rect 1851 479 1917 486
rect 1851 445 1867 479
rect 1901 445 1917 479
rect 1851 411 1917 445
rect 1851 377 1867 411
rect 1901 377 1917 411
rect 1851 343 1917 377
rect 1161 169 1287 203
rect 1127 153 1287 169
rect 564 55 586 89
rect 620 55 719 89
rect 753 89 793 105
rect 787 55 793 89
rect 841 73 861 107
rect 895 73 911 107
rect 945 73 961 107
rect 995 73 1093 107
rect 1143 101 1217 117
rect 395 17 461 55
rect 753 17 793 55
rect 1143 67 1177 101
rect 1211 67 1217 101
rect 1253 107 1287 153
rect 1321 191 1431 207
rect 1321 187 1367 191
rect 1321 153 1328 187
rect 1362 157 1367 187
rect 1401 157 1431 191
rect 1362 153 1431 157
rect 1321 141 1431 153
rect 1465 265 1525 281
rect 1708 265 1745 315
rect 1851 309 1867 343
rect 1901 309 1917 343
rect 1953 485 1987 527
rect 2143 485 2204 527
rect 1953 373 1987 451
rect 1953 323 1987 339
rect 2041 451 2057 485
rect 2091 451 2107 485
rect 2041 417 2107 451
rect 2041 383 2057 417
rect 2091 383 2107 417
rect 1851 306 1917 309
rect 1851 299 1923 306
rect 1882 286 1923 299
rect 1465 249 1674 265
rect 1465 215 1640 249
rect 1465 199 1674 215
rect 1708 249 1855 265
rect 1708 215 1821 249
rect 1708 199 1855 215
rect 1465 107 1499 199
rect 1708 165 1745 199
rect 1889 178 1923 286
rect 1882 165 1923 178
rect 1672 162 1745 165
rect 1672 128 1695 162
rect 1729 128 1745 162
rect 1851 158 1923 165
rect 2041 265 2107 383
rect 2143 451 2154 485
rect 2188 451 2204 485
rect 2322 485 2356 527
rect 2143 417 2204 451
rect 2143 383 2154 417
rect 2188 383 2204 417
rect 2143 349 2204 383
rect 2143 315 2154 349
rect 2188 315 2204 349
rect 2143 299 2204 315
rect 2238 449 2288 465
rect 2272 415 2288 449
rect 2238 381 2288 415
rect 2272 347 2288 381
rect 2238 289 2288 347
rect 2041 249 2213 265
rect 2041 215 2179 249
rect 2041 199 2213 215
rect 1851 157 1917 158
rect 1253 73 1295 107
rect 1329 73 1345 107
rect 1391 73 1407 107
rect 1441 73 1499 107
rect 1548 107 1622 123
rect 1548 73 1588 107
rect 1143 17 1217 67
rect 1548 17 1622 73
rect 1672 94 1745 128
rect 1672 60 1695 94
rect 1729 60 1745 94
rect 1779 123 1817 139
rect 1779 89 1781 123
rect 1815 89 1817 123
rect 1779 17 1817 89
rect 1851 123 1867 157
rect 1901 123 1917 157
rect 1851 89 1917 123
rect 1851 55 1867 89
rect 1901 55 1917 89
rect 1851 51 1917 55
rect 1951 122 1997 138
rect 1951 88 1953 122
rect 1987 88 1997 122
rect 1951 17 1997 88
rect 2041 119 2091 199
rect 2041 85 2057 119
rect 2041 69 2091 85
rect 2138 127 2154 161
rect 2188 127 2204 161
rect 2247 159 2288 289
rect 2322 417 2356 451
rect 2322 349 2356 383
rect 2322 279 2356 315
rect 2138 93 2204 127
rect 2138 59 2154 93
rect 2188 59 2204 93
rect 2138 17 2204 59
rect 2238 143 2288 159
rect 2272 109 2288 143
rect 2238 53 2288 109
rect 2322 161 2356 191
rect 2322 93 2356 127
rect 2322 17 2356 59
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 2053 527 2087 561
rect 2145 527 2179 561
rect 2237 527 2271 561
rect 2329 527 2363 561
rect 129 357 163 391
rect 210 153 244 187
rect 1041 365 1075 391
rect 1041 357 1045 365
rect 1045 357 1075 365
rect 949 153 983 187
rect 1325 357 1359 391
rect 1328 153 1362 187
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
rect 2053 -17 2087 17
rect 2145 -17 2179 17
rect 2237 -17 2271 17
rect 2329 -17 2363 17
<< metal1 >>
rect 0 561 2392 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2053 561
rect 2087 527 2145 561
rect 2179 527 2237 561
rect 2271 527 2329 561
rect 2363 527 2392 561
rect 0 496 2392 527
rect 117 391 175 397
rect 117 357 129 391
rect 163 388 175 391
rect 1029 391 1087 397
rect 1029 388 1041 391
rect 163 360 1041 388
rect 163 357 175 360
rect 117 351 175 357
rect 1029 357 1041 360
rect 1075 388 1087 391
rect 1313 391 1371 397
rect 1313 388 1325 391
rect 1075 360 1325 388
rect 1075 357 1087 360
rect 1029 351 1087 357
rect 1313 357 1325 360
rect 1359 357 1371 391
rect 1313 351 1371 357
rect 198 187 256 193
rect 198 153 210 187
rect 244 184 256 187
rect 937 187 995 193
rect 937 184 949 187
rect 244 156 949 184
rect 244 153 256 156
rect 198 147 256 153
rect 937 153 949 156
rect 983 184 995 187
rect 1316 187 1374 193
rect 1316 184 1328 187
rect 983 156 1328 184
rect 983 153 995 156
rect 937 147 995 153
rect 1316 153 1328 156
rect 1362 153 1374 187
rect 1316 147 1374 153
rect 0 17 2392 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2053 17
rect 2087 -17 2145 17
rect 2179 -17 2237 17
rect 2271 -17 2329 17
rect 2363 -17 2392 17
rect 0 -48 2392 -17
<< labels >>
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
flabel locali s 771 221 805 255 0 FreeSans 300 0 0 0 SCD
port 3 nsew signal input
flabel locali s 495 289 529 323 0 FreeSans 300 0 0 0 D
port 2 nsew signal input
flabel locali s 2247 289 2281 323 0 FreeSans 400 0 0 0 Q_N
port 10 nsew signal output
flabel locali s 495 85 529 119 0 FreeSans 300 0 0 0 SCE
port 4 nsew signal input
flabel locali s 31 221 65 255 0 FreeSans 400 0 0 0 CLK
port 1 nsew clock input
flabel locali s 1879 85 1913 119 0 FreeSans 200 0 0 0 Q
port 9 nsew signal output
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel pwell s 46 0 46 0 0 FreeSans 200 0 0 0 VNB
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel nwell s 46 544 46 544 0 FreeSans 200 0 0 0 VPB
rlabel comment s 0 0 0 0 4 sdfxbp_2
rlabel metal1 s 0 -48 2392 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2392 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2392 544
string GDS_END 361040
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 343158
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 11.960 0.000 
<< end >>
