magic
tech sky130A
magscale 1 2
timestamp 1704896540
<< nwell >>
rect -38 261 2062 582
<< pwell >>
rect 1 21 2023 203
rect 29 -17 63 21
<< scnmos >>
rect 79 47 109 177
rect 163 47 193 177
rect 484 47 514 177
rect 568 47 598 177
rect 652 47 682 177
rect 736 47 766 177
rect 820 47 850 177
rect 904 47 934 177
rect 988 47 1018 177
rect 1072 47 1102 177
rect 1324 47 1354 177
rect 1408 47 1438 177
rect 1492 47 1522 177
rect 1576 47 1606 177
rect 1660 47 1690 177
rect 1744 47 1774 177
rect 1828 47 1858 177
rect 1912 47 1942 177
<< scpmoshvt >>
rect 79 297 109 497
rect 163 297 193 497
rect 484 297 514 497
rect 568 297 598 497
rect 652 297 682 497
rect 736 297 766 497
rect 820 297 850 497
rect 904 297 934 497
rect 988 297 1018 497
rect 1072 297 1102 497
rect 1324 297 1354 497
rect 1408 297 1438 497
rect 1492 297 1522 497
rect 1576 297 1606 497
rect 1660 297 1690 497
rect 1744 297 1774 497
rect 1828 297 1858 497
rect 1912 297 1942 497
<< ndiff >>
rect 27 109 79 177
rect 27 75 35 109
rect 69 75 79 109
rect 27 47 79 75
rect 109 93 163 177
rect 109 59 119 93
rect 153 59 163 93
rect 109 47 163 59
rect 193 93 292 177
rect 193 59 219 93
rect 253 59 292 93
rect 193 47 292 59
rect 432 165 484 177
rect 432 131 440 165
rect 474 131 484 165
rect 432 47 484 131
rect 514 165 568 177
rect 514 131 524 165
rect 558 131 568 165
rect 514 47 568 131
rect 598 97 652 177
rect 598 63 608 97
rect 642 63 652 97
rect 598 47 652 63
rect 682 165 736 177
rect 682 131 692 165
rect 726 131 736 165
rect 682 47 736 131
rect 766 97 820 177
rect 766 63 776 97
rect 810 63 820 97
rect 766 47 820 63
rect 850 165 904 177
rect 850 131 860 165
rect 894 131 904 165
rect 850 47 904 131
rect 934 97 988 177
rect 934 63 944 97
rect 978 63 988 97
rect 934 47 988 63
rect 1018 165 1072 177
rect 1018 131 1028 165
rect 1062 131 1072 165
rect 1018 47 1072 131
rect 1102 97 1154 177
rect 1102 63 1112 97
rect 1146 63 1154 97
rect 1102 47 1154 63
rect 1266 165 1324 177
rect 1266 131 1280 165
rect 1314 131 1324 165
rect 1266 47 1324 131
rect 1354 97 1408 177
rect 1354 63 1364 97
rect 1398 63 1408 97
rect 1354 47 1408 63
rect 1438 165 1492 177
rect 1438 131 1448 165
rect 1482 131 1492 165
rect 1438 47 1492 131
rect 1522 97 1576 177
rect 1522 63 1532 97
rect 1566 63 1576 97
rect 1522 47 1576 63
rect 1606 165 1660 177
rect 1606 131 1616 165
rect 1650 131 1660 165
rect 1606 47 1660 131
rect 1690 97 1744 177
rect 1690 63 1700 97
rect 1734 63 1744 97
rect 1690 47 1744 63
rect 1774 165 1828 177
rect 1774 131 1784 165
rect 1818 131 1828 165
rect 1774 47 1828 131
rect 1858 97 1912 177
rect 1858 63 1868 97
rect 1902 63 1912 97
rect 1858 47 1912 63
rect 1942 165 1997 177
rect 1942 131 1952 165
rect 1986 131 1997 165
rect 1942 47 1997 131
<< pdiff >>
rect 27 472 79 497
rect 27 438 35 472
rect 69 438 79 472
rect 27 297 79 438
rect 109 489 163 497
rect 109 455 119 489
rect 153 455 163 489
rect 109 297 163 455
rect 193 483 292 497
rect 193 449 203 483
rect 237 449 292 483
rect 193 297 292 449
rect 432 485 484 497
rect 432 451 440 485
rect 474 451 484 485
rect 432 417 484 451
rect 432 383 440 417
rect 474 383 484 417
rect 432 349 484 383
rect 432 315 440 349
rect 474 315 484 349
rect 432 297 484 315
rect 514 477 568 497
rect 514 443 524 477
rect 558 443 568 477
rect 514 374 568 443
rect 514 340 524 374
rect 558 340 568 374
rect 514 297 568 340
rect 598 485 652 497
rect 598 451 608 485
rect 642 451 652 485
rect 598 417 652 451
rect 598 383 608 417
rect 642 383 652 417
rect 598 297 652 383
rect 682 485 736 497
rect 682 451 692 485
rect 726 451 736 485
rect 682 417 736 451
rect 682 383 692 417
rect 726 383 736 417
rect 682 349 736 383
rect 682 315 692 349
rect 726 315 736 349
rect 682 297 736 315
rect 766 485 820 497
rect 766 451 776 485
rect 810 451 820 485
rect 766 417 820 451
rect 766 383 776 417
rect 810 383 820 417
rect 766 297 820 383
rect 850 485 904 497
rect 850 451 860 485
rect 894 451 904 485
rect 850 417 904 451
rect 850 383 860 417
rect 894 383 904 417
rect 850 349 904 383
rect 850 315 860 349
rect 894 315 904 349
rect 850 297 904 315
rect 934 485 988 497
rect 934 451 944 485
rect 978 451 988 485
rect 934 417 988 451
rect 934 383 944 417
rect 978 383 988 417
rect 934 297 988 383
rect 1018 485 1072 497
rect 1018 451 1028 485
rect 1062 451 1072 485
rect 1018 417 1072 451
rect 1018 383 1028 417
rect 1062 383 1072 417
rect 1018 349 1072 383
rect 1018 315 1028 349
rect 1062 315 1072 349
rect 1018 297 1072 315
rect 1102 485 1324 497
rect 1102 451 1122 485
rect 1156 451 1191 485
rect 1225 451 1274 485
rect 1308 451 1324 485
rect 1102 417 1324 451
rect 1102 383 1122 417
rect 1156 383 1191 417
rect 1225 383 1274 417
rect 1308 383 1324 417
rect 1102 297 1324 383
rect 1354 485 1408 497
rect 1354 451 1364 485
rect 1398 451 1408 485
rect 1354 417 1408 451
rect 1354 383 1364 417
rect 1398 383 1408 417
rect 1354 349 1408 383
rect 1354 315 1364 349
rect 1398 315 1408 349
rect 1354 297 1408 315
rect 1438 485 1492 497
rect 1438 451 1448 485
rect 1482 451 1492 485
rect 1438 417 1492 451
rect 1438 383 1448 417
rect 1482 383 1492 417
rect 1438 297 1492 383
rect 1522 485 1576 497
rect 1522 451 1532 485
rect 1566 451 1576 485
rect 1522 417 1576 451
rect 1522 383 1532 417
rect 1566 383 1576 417
rect 1522 349 1576 383
rect 1522 315 1532 349
rect 1566 315 1576 349
rect 1522 297 1576 315
rect 1606 485 1660 497
rect 1606 451 1616 485
rect 1650 451 1660 485
rect 1606 417 1660 451
rect 1606 383 1616 417
rect 1650 383 1660 417
rect 1606 297 1660 383
rect 1690 485 1744 497
rect 1690 451 1700 485
rect 1734 451 1744 485
rect 1690 417 1744 451
rect 1690 383 1700 417
rect 1734 383 1744 417
rect 1690 349 1744 383
rect 1690 315 1700 349
rect 1734 315 1744 349
rect 1690 297 1744 315
rect 1774 485 1828 497
rect 1774 451 1784 485
rect 1818 451 1828 485
rect 1774 417 1828 451
rect 1774 383 1784 417
rect 1818 383 1828 417
rect 1774 297 1828 383
rect 1858 485 1912 497
rect 1858 451 1868 485
rect 1902 451 1912 485
rect 1858 417 1912 451
rect 1858 383 1868 417
rect 1902 383 1912 417
rect 1858 349 1912 383
rect 1858 315 1868 349
rect 1902 315 1912 349
rect 1858 297 1912 315
rect 1942 485 1997 497
rect 1942 451 1952 485
rect 1986 451 1997 485
rect 1942 417 1997 451
rect 1942 383 1952 417
rect 1986 383 1997 417
rect 1942 349 1997 383
rect 1942 315 1952 349
rect 1986 315 1997 349
rect 1942 297 1997 315
<< ndiffc >>
rect 35 75 69 109
rect 119 59 153 93
rect 219 59 253 93
rect 440 131 474 165
rect 524 131 558 165
rect 608 63 642 97
rect 692 131 726 165
rect 776 63 810 97
rect 860 131 894 165
rect 944 63 978 97
rect 1028 131 1062 165
rect 1112 63 1146 97
rect 1280 131 1314 165
rect 1364 63 1398 97
rect 1448 131 1482 165
rect 1532 63 1566 97
rect 1616 131 1650 165
rect 1700 63 1734 97
rect 1784 131 1818 165
rect 1868 63 1902 97
rect 1952 131 1986 165
<< pdiffc >>
rect 35 438 69 472
rect 119 455 153 489
rect 203 449 237 483
rect 440 451 474 485
rect 440 383 474 417
rect 440 315 474 349
rect 524 443 558 477
rect 524 340 558 374
rect 608 451 642 485
rect 608 383 642 417
rect 692 451 726 485
rect 692 383 726 417
rect 692 315 726 349
rect 776 451 810 485
rect 776 383 810 417
rect 860 451 894 485
rect 860 383 894 417
rect 860 315 894 349
rect 944 451 978 485
rect 944 383 978 417
rect 1028 451 1062 485
rect 1028 383 1062 417
rect 1028 315 1062 349
rect 1122 451 1156 485
rect 1191 451 1225 485
rect 1274 451 1308 485
rect 1122 383 1156 417
rect 1191 383 1225 417
rect 1274 383 1308 417
rect 1364 451 1398 485
rect 1364 383 1398 417
rect 1364 315 1398 349
rect 1448 451 1482 485
rect 1448 383 1482 417
rect 1532 451 1566 485
rect 1532 383 1566 417
rect 1532 315 1566 349
rect 1616 451 1650 485
rect 1616 383 1650 417
rect 1700 451 1734 485
rect 1700 383 1734 417
rect 1700 315 1734 349
rect 1784 451 1818 485
rect 1784 383 1818 417
rect 1868 451 1902 485
rect 1868 383 1902 417
rect 1868 315 1902 349
rect 1952 451 1986 485
rect 1952 383 1986 417
rect 1952 315 1986 349
<< poly >>
rect 79 497 109 523
rect 163 497 193 523
rect 484 497 514 523
rect 568 497 598 523
rect 652 497 682 523
rect 736 497 766 523
rect 820 497 850 523
rect 904 497 934 523
rect 988 497 1018 523
rect 1072 497 1102 523
rect 1324 497 1354 523
rect 1408 497 1438 523
rect 1492 497 1522 523
rect 1576 497 1606 523
rect 1660 497 1690 523
rect 1744 497 1774 523
rect 1828 497 1858 523
rect 1912 497 1942 523
rect 79 265 109 297
rect 163 265 193 297
rect 484 265 514 297
rect 21 249 109 265
rect 21 215 32 249
rect 66 215 109 249
rect 21 199 109 215
rect 151 249 205 265
rect 151 215 161 249
rect 195 215 205 249
rect 151 199 205 215
rect 247 259 514 265
rect 568 259 598 297
rect 652 259 682 297
rect 736 259 766 297
rect 247 249 766 259
rect 247 215 257 249
rect 291 215 524 249
rect 558 215 607 249
rect 641 215 766 249
rect 247 205 766 215
rect 247 199 514 205
rect 79 177 109 199
rect 163 177 193 199
rect 484 177 514 199
rect 568 177 598 205
rect 652 177 682 205
rect 736 177 766 205
rect 820 259 850 297
rect 904 259 934 297
rect 988 259 1018 297
rect 1072 259 1102 297
rect 1324 259 1354 297
rect 1408 259 1438 297
rect 1492 259 1522 297
rect 1576 259 1606 297
rect 820 249 1102 259
rect 820 215 861 249
rect 895 215 943 249
rect 977 215 1028 249
rect 1062 215 1102 249
rect 820 205 1102 215
rect 1258 249 1606 259
rect 1258 215 1274 249
rect 1308 215 1364 249
rect 1398 215 1448 249
rect 1482 215 1532 249
rect 1566 215 1606 249
rect 1258 205 1606 215
rect 820 177 850 205
rect 904 177 934 205
rect 988 177 1018 205
rect 1072 177 1102 205
rect 1324 177 1354 205
rect 1408 177 1438 205
rect 1492 177 1522 205
rect 1576 177 1606 205
rect 1660 259 1690 297
rect 1744 259 1774 297
rect 1828 259 1858 297
rect 1912 261 1942 297
rect 1912 259 2003 261
rect 1660 249 2003 259
rect 1660 215 1700 249
rect 1734 215 1784 249
rect 1818 215 1868 249
rect 1902 215 1952 249
rect 1986 215 2003 249
rect 1660 205 2003 215
rect 1660 177 1690 205
rect 1744 177 1774 205
rect 1828 177 1858 205
rect 1912 203 2003 205
rect 1912 177 1942 203
rect 79 21 109 47
rect 163 21 193 47
rect 484 21 514 47
rect 568 21 598 47
rect 652 21 682 47
rect 736 21 766 47
rect 820 21 850 47
rect 904 21 934 47
rect 988 21 1018 47
rect 1072 21 1102 47
rect 1324 21 1354 47
rect 1408 21 1438 47
rect 1492 21 1522 47
rect 1576 21 1606 47
rect 1660 21 1690 47
rect 1744 21 1774 47
rect 1828 21 1858 47
rect 1912 21 1942 47
<< polycont >>
rect 32 215 66 249
rect 161 215 195 249
rect 257 215 291 249
rect 524 215 558 249
rect 607 215 641 249
rect 861 215 895 249
rect 943 215 977 249
rect 1028 215 1062 249
rect 1274 215 1308 249
rect 1364 215 1398 249
rect 1448 215 1482 249
rect 1532 215 1566 249
rect 1700 215 1734 249
rect 1784 215 1818 249
rect 1868 215 1902 249
rect 1952 215 1986 249
<< locali >>
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 108 489 153 527
rect 17 472 74 488
rect 17 438 35 472
rect 69 438 74 472
rect 108 455 119 489
rect 108 439 153 455
rect 187 483 359 493
rect 187 449 203 483
rect 237 449 359 483
rect 17 396 74 438
rect 187 430 359 449
rect 17 357 291 396
rect 20 249 66 323
rect 20 215 32 249
rect 20 199 66 215
rect 118 249 195 323
rect 118 215 161 249
rect 118 199 195 215
rect 229 249 291 357
rect 229 215 257 249
rect 229 161 291 215
rect 17 127 291 161
rect 325 261 359 430
rect 440 485 474 527
rect 440 417 474 451
rect 440 349 474 383
rect 440 299 474 315
rect 508 477 558 493
rect 508 443 524 477
rect 508 374 558 443
rect 508 340 524 374
rect 592 485 642 527
rect 592 451 608 485
rect 592 417 642 451
rect 592 383 608 417
rect 592 367 642 383
rect 676 485 742 493
rect 676 451 692 485
rect 726 451 742 485
rect 676 417 742 451
rect 676 383 692 417
rect 726 383 742 417
rect 508 333 558 340
rect 676 349 742 383
rect 776 485 810 527
rect 776 417 810 451
rect 776 367 810 383
rect 844 485 910 493
rect 844 451 860 485
rect 894 451 910 485
rect 844 417 910 451
rect 844 383 860 417
rect 894 383 910 417
rect 676 333 692 349
rect 508 315 692 333
rect 726 333 742 349
rect 844 349 910 383
rect 944 485 978 527
rect 944 417 978 451
rect 944 367 978 383
rect 1012 485 1078 493
rect 1012 451 1028 485
rect 1062 451 1078 485
rect 1012 417 1078 451
rect 1012 383 1028 417
rect 1062 383 1078 417
rect 844 333 860 349
rect 726 315 860 333
rect 894 333 910 349
rect 1012 349 1078 383
rect 1122 485 1308 527
rect 1156 451 1191 485
rect 1225 451 1274 485
rect 1122 417 1308 451
rect 1156 383 1191 417
rect 1225 383 1274 417
rect 1122 367 1308 383
rect 1348 485 1414 493
rect 1348 451 1364 485
rect 1398 451 1414 485
rect 1348 417 1414 451
rect 1348 383 1364 417
rect 1398 383 1414 417
rect 1012 333 1028 349
rect 894 315 1028 333
rect 1062 333 1078 349
rect 1348 349 1414 383
rect 1448 485 1482 527
rect 1448 417 1482 451
rect 1448 367 1482 383
rect 1516 485 1582 493
rect 1516 451 1532 485
rect 1566 451 1582 485
rect 1516 417 1582 451
rect 1516 383 1532 417
rect 1566 383 1582 417
rect 1348 333 1364 349
rect 1062 315 1364 333
rect 1398 333 1414 349
rect 1516 349 1582 383
rect 1616 485 1650 527
rect 1616 417 1650 451
rect 1616 367 1650 383
rect 1684 485 1750 493
rect 1684 451 1700 485
rect 1734 451 1750 485
rect 1684 417 1750 451
rect 1684 383 1700 417
rect 1734 383 1750 417
rect 1516 333 1532 349
rect 1398 315 1532 333
rect 1566 333 1582 349
rect 1684 349 1750 383
rect 1784 485 1818 527
rect 1784 417 1818 451
rect 1784 367 1818 383
rect 1852 485 1918 493
rect 1852 451 1868 485
rect 1902 451 1918 485
rect 1852 417 1918 451
rect 1852 383 1868 417
rect 1902 383 1918 417
rect 1684 333 1700 349
rect 1566 315 1700 333
rect 1734 333 1750 349
rect 1852 349 1918 383
rect 1852 333 1868 349
rect 1734 315 1868 333
rect 1902 315 1918 349
rect 508 289 1918 315
rect 1952 485 2007 527
rect 1986 451 2007 485
rect 1952 417 2007 451
rect 1986 383 2007 417
rect 1952 349 2007 383
rect 1986 315 2007 349
rect 1952 289 2007 315
rect 325 255 442 261
rect 325 221 396 255
rect 430 221 442 255
rect 325 215 442 221
rect 508 215 524 249
rect 558 215 607 249
rect 641 215 657 249
rect 17 109 69 127
rect 17 75 35 109
rect 325 93 359 215
rect 740 181 798 289
rect 832 221 856 255
rect 890 249 1078 255
rect 832 215 861 221
rect 895 215 943 249
rect 977 215 1028 249
rect 1062 215 1078 249
rect 1224 249 1582 255
rect 1224 215 1274 249
rect 1308 215 1364 249
rect 1398 215 1448 249
rect 1482 215 1532 249
rect 1566 215 1582 249
rect 1684 249 2003 255
rect 1684 215 1700 249
rect 1734 215 1784 249
rect 1818 215 1868 249
rect 1902 215 1952 249
rect 1986 215 2003 249
rect 17 51 69 75
rect 103 59 119 93
rect 153 59 169 93
rect 103 17 169 59
rect 203 59 219 93
rect 253 59 359 93
rect 203 51 359 59
rect 440 165 474 181
rect 508 165 798 181
rect 508 131 524 165
rect 558 131 692 165
rect 726 131 798 165
rect 844 165 1230 181
rect 844 131 860 165
rect 894 131 1028 165
rect 1062 147 1230 165
rect 1062 131 1078 147
rect 440 97 474 131
rect 1196 97 1230 147
rect 1264 165 2007 181
rect 1264 131 1280 165
rect 1314 131 1448 165
rect 1482 131 1616 165
rect 1650 131 1784 165
rect 1818 131 1952 165
rect 1986 131 2007 165
rect 440 63 608 97
rect 642 63 776 97
rect 810 63 944 97
rect 978 63 1112 97
rect 1146 63 1162 97
rect 440 51 1162 63
rect 1196 63 1364 97
rect 1398 63 1532 97
rect 1566 63 1582 97
rect 1196 51 1582 63
rect 1684 63 1700 97
rect 1734 63 1750 97
rect 1684 17 1750 63
rect 1852 63 1868 97
rect 1902 63 1918 97
rect 1852 17 1918 63
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
<< viali >>
rect 29 527 63 561
rect 121 527 155 561
rect 213 527 247 561
rect 305 527 339 561
rect 397 527 431 561
rect 489 527 523 561
rect 581 527 615 561
rect 673 527 707 561
rect 765 527 799 561
rect 857 527 891 561
rect 949 527 983 561
rect 1041 527 1075 561
rect 1133 527 1167 561
rect 1225 527 1259 561
rect 1317 527 1351 561
rect 1409 527 1443 561
rect 1501 527 1535 561
rect 1593 527 1627 561
rect 1685 527 1719 561
rect 1777 527 1811 561
rect 1869 527 1903 561
rect 1961 527 1995 561
rect 396 221 430 255
rect 856 249 890 255
rect 856 221 861 249
rect 861 221 890 249
rect 29 -17 63 17
rect 121 -17 155 17
rect 213 -17 247 17
rect 305 -17 339 17
rect 397 -17 431 17
rect 489 -17 523 17
rect 581 -17 615 17
rect 673 -17 707 17
rect 765 -17 799 17
rect 857 -17 891 17
rect 949 -17 983 17
rect 1041 -17 1075 17
rect 1133 -17 1167 17
rect 1225 -17 1259 17
rect 1317 -17 1351 17
rect 1409 -17 1443 17
rect 1501 -17 1535 17
rect 1593 -17 1627 17
rect 1685 -17 1719 17
rect 1777 -17 1811 17
rect 1869 -17 1903 17
rect 1961 -17 1995 17
<< metal1 >>
rect 0 561 2024 592
rect 0 527 29 561
rect 63 527 121 561
rect 155 527 213 561
rect 247 527 305 561
rect 339 527 397 561
rect 431 527 489 561
rect 523 527 581 561
rect 615 527 673 561
rect 707 527 765 561
rect 799 527 857 561
rect 891 527 949 561
rect 983 527 1041 561
rect 1075 527 1133 561
rect 1167 527 1225 561
rect 1259 527 1317 561
rect 1351 527 1409 561
rect 1443 527 1501 561
rect 1535 527 1593 561
rect 1627 527 1685 561
rect 1719 527 1777 561
rect 1811 527 1869 561
rect 1903 527 1961 561
rect 1995 527 2024 561
rect 0 496 2024 527
rect 384 255 442 261
rect 384 221 396 255
rect 430 252 442 255
rect 844 255 902 261
rect 844 252 856 255
rect 430 224 856 252
rect 430 221 442 224
rect 384 215 442 221
rect 844 221 856 224
rect 890 221 902 255
rect 844 215 902 221
rect 0 17 2024 48
rect 0 -17 29 17
rect 63 -17 121 17
rect 155 -17 213 17
rect 247 -17 305 17
rect 339 -17 397 17
rect 431 -17 489 17
rect 523 -17 581 17
rect 615 -17 673 17
rect 707 -17 765 17
rect 799 -17 857 17
rect 891 -17 949 17
rect 983 -17 1041 17
rect 1075 -17 1133 17
rect 1167 -17 1225 17
rect 1259 -17 1317 17
rect 1351 -17 1409 17
rect 1443 -17 1501 17
rect 1535 -17 1593 17
rect 1627 -17 1685 17
rect 1719 -17 1777 17
rect 1811 -17 1869 17
rect 1903 -17 1961 17
rect 1995 -17 2024 17
rect 0 -48 2024 -17
<< labels >>
flabel locali s 122 221 156 255 0 FreeSans 200 0 0 0 B_N
port 2 nsew signal input
flabel locali s 30 221 64 255 0 FreeSans 200 0 0 0 A_N
port 1 nsew signal input
flabel locali s 1224 221 1258 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 764 153 798 187 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 764 289 798 323 0 FreeSans 200 0 0 0 Y
port 9 nsew signal output
flabel locali s 1316 221 1350 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1408 221 1442 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1500 221 1534 255 0 FreeSans 200 0 0 0 C
port 3 nsew signal input
flabel locali s 1684 221 1718 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 1868 221 1902 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 1960 221 1994 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel locali s 1776 221 1810 255 0 FreeSans 200 0 0 0 D
port 4 nsew signal input
flabel pwell s 29 -17 63 17 0 FreeSans 200 0 0 0 VNB
port 6 nsew ground bidirectional
flabel nwell s 29 527 63 561 0 FreeSans 200 0 0 0 VPB
port 7 nsew power bidirectional
flabel metal1 s 29 -17 63 17 0 FreeSans 200 0 0 0 VGND
port 5 nsew ground bidirectional abutment
flabel metal1 s 29 527 63 561 0 FreeSans 200 0 0 0 VPWR
port 8 nsew power bidirectional abutment
rlabel comment s 0 0 0 0 4 nand4bb_4
rlabel metal1 s 0 -48 2024 48 1 VGND
port 5 nsew ground bidirectional abutment
rlabel metal1 s 0 496 2024 592 1 VPWR
port 8 nsew power bidirectional abutment
<< properties >>
string FIXED_BBOX 0 0 2024 544
string GDS_END 1953980
string GDS_FILE $PDKPATH/libs.ref/sky130_fd_sc_hd/gds/sky130_fd_sc_hd.gds
string GDS_START 1938992
string LEFclass CORE
string LEFsite unithd
string LEFsymmetry X Y R90
string path 0.000 0.000 50.600 0.000 
<< end >>
